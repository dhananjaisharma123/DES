
--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_in_pkg_v1 IS

COMPONENT ccs_in_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    idat   : OUT std_logic_vector(width-1 DOWNTO 0);
    dat    : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_in_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_in_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    idat  : OUT std_logic_vector(width-1 DOWNTO 0);
    dat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_in_v1;

ARCHITECTURE beh OF ccs_in_v1 IS
BEGIN

  idat <= dat;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_out_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_out_pkg_v1 IS

COMPONENT ccs_out_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    dat    : OUT std_logic_vector(width-1 DOWNTO 0);
    idat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_out_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_out_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    dat   : OUT std_logic_vector(width-1 DOWNTO 0);
    idat  : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_out_v1;

ARCHITECTURE beh OF ccs_out_v1 IS
BEGIN

  dat <= idat;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_io_sync_pkg_v2 IS

COMPONENT mgc_io_sync_v2
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END COMPONENT;

END mgc_io_sync_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_io_sync_v2 IS
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END mgc_io_sync_v2;

ARCHITECTURE beh OF mgc_io_sync_v2 IS
BEGIN

  lz <= ld;

END beh;


--------> ./rtl_des_checkmgc_rom_12_512_4_1.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   ds6365@hansolo.poly.edu
--  Generated date: Sun Mar 21 12:47:51 2021
-- ----------------------------------------------------------------------

-- 
LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


PACKAGE des_checkmgc_rom_12_512_4_1_pkg IS 
  COMPONENT des_checkmgc_rom_12_512_4_1
    PORT (
      addr : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
      data_out : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
  END COMPONENT;
END des_checkmgc_rom_12_512_4_1_pkg;

PACKAGE BODY des_checkmgc_rom_12_512_4_1_pkg IS
END des_checkmgc_rom_12_512_4_1_pkg;

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


USE work.des_checkmgc_rom_12_512_4_1_pkg.all;
LIBRARY std;

USE std.textio.all;
USE ieee.std_logic_textio.all;

ENTITY des_checkmgc_rom_12_512_4_1 IS
    PORT (
      addr : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
      data_out : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END des_checkmgc_rom_12_512_4_1;

ARCHITECTURE v1 OF des_checkmgc_rom_12_512_4_1 IS
  -- Start of SIF_NL_VHDL::nhl_rom_body
  -- Constants for ROM dimensions
  CONSTANT n_width    : INTEGER := 4;
  CONSTANT n_size     : INTEGER := 512;
  CONSTANT n_addr_w   : INTEGER := 9;
  CONSTANT n_inreg    : INTEGER := 0;
  CONSTANT n_outreg   : INTEGER := 0;
  -- Define data types for ROM storage;
  SUBTYPE  word  IS std_logic_vector((n_width)-1 DOWNTO 0);
  TYPE     table IS ARRAY (0 to n_size-1) of word;

  SIGNAL mem : table := table'(
    word'("1110"),
    word'("0100"),
    word'("1101"),
    word'("0001"),
    word'("0010"),
    word'("1111"),
    word'("1011"),
    word'("1000"),
    word'("0011"),
    word'("1010"),
    word'("0110"),
    word'("1100"),
    word'("0101"),
    word'("1001"),
    word'("0000"),
    word'("0111"),
    word'("0000"),
    word'("1111"),
    word'("0111"),
    word'("0100"),
    word'("1110"),
    word'("0010"),
    word'("1101"),
    word'("0001"),
    word'("1010"),
    word'("0110"),
    word'("1100"),
    word'("1011"),
    word'("1001"),
    word'("0101"),
    word'("0011"),
    word'("1000"),
    word'("0100"),
    word'("0001"),
    word'("1110"),
    word'("1000"),
    word'("1101"),
    word'("0110"),
    word'("0010"),
    word'("1011"),
    word'("1111"),
    word'("1100"),
    word'("1001"),
    word'("0111"),
    word'("0011"),
    word'("1010"),
    word'("0101"),
    word'("0000"),
    word'("1111"),
    word'("1100"),
    word'("1000"),
    word'("0010"),
    word'("0100"),
    word'("1001"),
    word'("0001"),
    word'("0111"),
    word'("0101"),
    word'("1011"),
    word'("0011"),
    word'("1110"),
    word'("1010"),
    word'("0000"),
    word'("0110"),
    word'("1101"),
    word'("1111"),
    word'("0001"),
    word'("1000"),
    word'("1110"),
    word'("0110"),
    word'("1011"),
    word'("0011"),
    word'("0100"),
    word'("1001"),
    word'("0111"),
    word'("0010"),
    word'("1101"),
    word'("1100"),
    word'("0000"),
    word'("0101"),
    word'("1010"),
    word'("0011"),
    word'("1101"),
    word'("0100"),
    word'("0111"),
    word'("1111"),
    word'("0010"),
    word'("1000"),
    word'("1110"),
    word'("1100"),
    word'("0000"),
    word'("0001"),
    word'("1010"),
    word'("0110"),
    word'("1001"),
    word'("1011"),
    word'("0101"),
    word'("0000"),
    word'("1110"),
    word'("0111"),
    word'("1011"),
    word'("1010"),
    word'("0100"),
    word'("1101"),
    word'("0001"),
    word'("0101"),
    word'("1000"),
    word'("1100"),
    word'("0110"),
    word'("1001"),
    word'("0011"),
    word'("0010"),
    word'("1111"),
    word'("1101"),
    word'("1000"),
    word'("1010"),
    word'("0001"),
    word'("0011"),
    word'("1111"),
    word'("0100"),
    word'("0010"),
    word'("1011"),
    word'("0110"),
    word'("0111"),
    word'("1100"),
    word'("0000"),
    word'("0101"),
    word'("1110"),
    word'("1001"),
    word'("1010"),
    word'("0000"),
    word'("1001"),
    word'("1110"),
    word'("0110"),
    word'("0011"),
    word'("1111"),
    word'("0101"),
    word'("0001"),
    word'("1101"),
    word'("1100"),
    word'("0111"),
    word'("1011"),
    word'("0100"),
    word'("0010"),
    word'("1000"),
    word'("1101"),
    word'("0111"),
    word'("0000"),
    word'("1001"),
    word'("0011"),
    word'("0100"),
    word'("0110"),
    word'("1010"),
    word'("0010"),
    word'("1000"),
    word'("0101"),
    word'("1110"),
    word'("1100"),
    word'("1011"),
    word'("1111"),
    word'("0001"),
    word'("1101"),
    word'("0110"),
    word'("0100"),
    word'("1001"),
    word'("1000"),
    word'("1111"),
    word'("0011"),
    word'("0000"),
    word'("1011"),
    word'("0001"),
    word'("0010"),
    word'("1100"),
    word'("0101"),
    word'("1010"),
    word'("1110"),
    word'("0111"),
    word'("0001"),
    word'("1010"),
    word'("1101"),
    word'("0000"),
    word'("0110"),
    word'("1001"),
    word'("1000"),
    word'("0111"),
    word'("0100"),
    word'("1111"),
    word'("1110"),
    word'("0011"),
    word'("1011"),
    word'("0101"),
    word'("0010"),
    word'("1100"),
    word'("0111"),
    word'("1101"),
    word'("1110"),
    word'("0011"),
    word'("0000"),
    word'("0110"),
    word'("1001"),
    word'("1010"),
    word'("0001"),
    word'("0010"),
    word'("1000"),
    word'("0101"),
    word'("1011"),
    word'("1100"),
    word'("0100"),
    word'("1111"),
    word'("1101"),
    word'("1000"),
    word'("1011"),
    word'("0101"),
    word'("0110"),
    word'("1111"),
    word'("0000"),
    word'("0011"),
    word'("0100"),
    word'("0111"),
    word'("0010"),
    word'("1100"),
    word'("0001"),
    word'("1010"),
    word'("1110"),
    word'("1001"),
    word'("1010"),
    word'("0110"),
    word'("1001"),
    word'("0000"),
    word'("1100"),
    word'("1011"),
    word'("0111"),
    word'("1101"),
    word'("1111"),
    word'("0001"),
    word'("0011"),
    word'("1110"),
    word'("0101"),
    word'("0010"),
    word'("1000"),
    word'("0100"),
    word'("0011"),
    word'("1111"),
    word'("0000"),
    word'("0110"),
    word'("1010"),
    word'("0001"),
    word'("1101"),
    word'("1000"),
    word'("1001"),
    word'("0100"),
    word'("0101"),
    word'("1011"),
    word'("1100"),
    word'("0111"),
    word'("0010"),
    word'("1110"),
    word'("0010"),
    word'("1100"),
    word'("0100"),
    word'("0001"),
    word'("0111"),
    word'("1010"),
    word'("1011"),
    word'("0110"),
    word'("1000"),
    word'("0101"),
    word'("0011"),
    word'("1111"),
    word'("1101"),
    word'("0000"),
    word'("1110"),
    word'("1001"),
    word'("1110"),
    word'("1011"),
    word'("0010"),
    word'("1100"),
    word'("0100"),
    word'("0111"),
    word'("1101"),
    word'("0001"),
    word'("0101"),
    word'("0000"),
    word'("1111"),
    word'("1010"),
    word'("0011"),
    word'("1001"),
    word'("1000"),
    word'("0110"),
    word'("0100"),
    word'("0010"),
    word'("0001"),
    word'("1011"),
    word'("1010"),
    word'("1101"),
    word'("0111"),
    word'("1000"),
    word'("1111"),
    word'("1001"),
    word'("1100"),
    word'("0101"),
    word'("0110"),
    word'("0011"),
    word'("0000"),
    word'("1110"),
    word'("1011"),
    word'("1000"),
    word'("1100"),
    word'("0111"),
    word'("0001"),
    word'("1110"),
    word'("0010"),
    word'("1101"),
    word'("0110"),
    word'("1111"),
    word'("0000"),
    word'("1001"),
    word'("1010"),
    word'("0100"),
    word'("0101"),
    word'("0011"),
    word'("1100"),
    word'("0001"),
    word'("1010"),
    word'("1111"),
    word'("1001"),
    word'("0010"),
    word'("0110"),
    word'("1000"),
    word'("0000"),
    word'("1101"),
    word'("0011"),
    word'("0100"),
    word'("1110"),
    word'("0111"),
    word'("0101"),
    word'("1011"),
    word'("1010"),
    word'("1111"),
    word'("0100"),
    word'("0010"),
    word'("0111"),
    word'("1100"),
    word'("1001"),
    word'("0101"),
    word'("0110"),
    word'("0001"),
    word'("1101"),
    word'("1110"),
    word'("0000"),
    word'("1011"),
    word'("0011"),
    word'("1000"),
    word'("1001"),
    word'("1110"),
    word'("1111"),
    word'("0101"),
    word'("0010"),
    word'("1000"),
    word'("1100"),
    word'("0011"),
    word'("0111"),
    word'("0000"),
    word'("0100"),
    word'("1010"),
    word'("0001"),
    word'("1101"),
    word'("1011"),
    word'("0110"),
    word'("0100"),
    word'("0011"),
    word'("0010"),
    word'("1100"),
    word'("1001"),
    word'("0101"),
    word'("1111"),
    word'("1010"),
    word'("1011"),
    word'("1110"),
    word'("0001"),
    word'("0111"),
    word'("0110"),
    word'("0000"),
    word'("1000"),
    word'("1101"),
    word'("0100"),
    word'("1011"),
    word'("0010"),
    word'("1110"),
    word'("1111"),
    word'("0000"),
    word'("1000"),
    word'("1101"),
    word'("0011"),
    word'("1100"),
    word'("1001"),
    word'("0111"),
    word'("0101"),
    word'("1010"),
    word'("0110"),
    word'("0001"),
    word'("1101"),
    word'("0000"),
    word'("1011"),
    word'("0111"),
    word'("0100"),
    word'("1001"),
    word'("0001"),
    word'("1010"),
    word'("1110"),
    word'("0011"),
    word'("0101"),
    word'("1100"),
    word'("0010"),
    word'("1111"),
    word'("1000"),
    word'("0110"),
    word'("0001"),
    word'("0100"),
    word'("1011"),
    word'("1101"),
    word'("1100"),
    word'("0011"),
    word'("0111"),
    word'("1110"),
    word'("1010"),
    word'("1111"),
    word'("0110"),
    word'("1000"),
    word'("0000"),
    word'("0101"),
    word'("1001"),
    word'("0010"),
    word'("0110"),
    word'("1011"),
    word'("1101"),
    word'("1000"),
    word'("0001"),
    word'("0100"),
    word'("1010"),
    word'("0111"),
    word'("1001"),
    word'("0101"),
    word'("0000"),
    word'("1111"),
    word'("1110"),
    word'("0010"),
    word'("0011"),
    word'("1100"),
    word'("1101"),
    word'("0010"),
    word'("1000"),
    word'("0100"),
    word'("0110"),
    word'("1111"),
    word'("1011"),
    word'("0001"),
    word'("1010"),
    word'("1001"),
    word'("0011"),
    word'("1110"),
    word'("0101"),
    word'("0000"),
    word'("1100"),
    word'("0111"),
    word'("0001"),
    word'("1111"),
    word'("1101"),
    word'("1000"),
    word'("1010"),
    word'("0011"),
    word'("0111"),
    word'("0100"),
    word'("1100"),
    word'("0101"),
    word'("0110"),
    word'("1011"),
    word'("0000"),
    word'("1110"),
    word'("1001"),
    word'("0010"),
    word'("0111"),
    word'("1011"),
    word'("0100"),
    word'("0001"),
    word'("1001"),
    word'("1100"),
    word'("1110"),
    word'("0010"),
    word'("0000"),
    word'("0110"),
    word'("1010"),
    word'("1101"),
    word'("1111"),
    word'("0011"),
    word'("0101"),
    word'("1000"),
    word'("0010"),
    word'("0001"),
    word'("1110"),
    word'("0111"),
    word'("0100"),
    word'("1010"),
    word'("1000"),
    word'("1101"),
    word'("1111"),
    word'("1100"),
    word'("1001"),
    word'("0000"),
    word'("0011"),
    word'("0101"),
    word'("0110"),
    word'("1011")
  );
  ATTRIBUTE rom_style : string;
  ATTRIBUTE rom_style OF mem : SIGNAL IS "block";
BEGIN

  -- Reading ROM
  PROCESS(addr)
    VARIABLE idx_addr : INTEGER;
  BEGIN
    idx_addr := conv_integer(unsigned(addr(8 DOWNTO 0)));
    data_out <= mem(idx_addr);
  END PROCESS;

END v1;



--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   ds6365@hansolo.poly.edu
--  Generated date: Sun Mar 21 12:47:50 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    des_check_core_core_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;


ENTITY des_check_core_core_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (16 DOWNTO 0)
  );
END des_check_core_core_fsm;

ARCHITECTURE v1 OF des_check_core_core_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for des_check_core_core_fsm_1
  TYPE des_check_core_core_fsm_1_ST IS (main_C_0, main_C_1, main_C_2, main_C_3, main_C_4,
      main_C_5, main_C_6, main_C_7, main_C_8, main_C_9, main_C_10, main_C_11, main_C_12,
      main_C_13, main_C_14, main_C_15, main_C_16);

  SIGNAL state_var : des_check_core_core_fsm_1_ST;
  SIGNAL state_var_NS : des_check_core_core_fsm_1_ST;

BEGIN
  des_check_core_core_fsm_1 : PROCESS (state_var)
  BEGIN
    CASE state_var IS
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000010");
        state_var_NS <= main_C_2;
      WHEN main_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000100");
        state_var_NS <= main_C_3;
      WHEN main_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000001000");
        state_var_NS <= main_C_4;
      WHEN main_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000010000");
        state_var_NS <= main_C_5;
      WHEN main_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000100000");
        state_var_NS <= main_C_6;
      WHEN main_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000001000000");
        state_var_NS <= main_C_7;
      WHEN main_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000010000000");
        state_var_NS <= main_C_8;
      WHEN main_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000100000000");
        state_var_NS <= main_C_9;
      WHEN main_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001000000000");
        state_var_NS <= main_C_10;
      WHEN main_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010000000000");
        state_var_NS <= main_C_11;
      WHEN main_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100000000000");
        state_var_NS <= main_C_12;
      WHEN main_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000000000000");
        state_var_NS <= main_C_13;
      WHEN main_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000000000000");
        state_var_NS <= main_C_14;
      WHEN main_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000000000000");
        state_var_NS <= main_C_15;
      WHEN main_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000000000000");
        state_var_NS <= main_C_16;
      WHEN main_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000000000000");
        state_var_NS <= main_C_0;
      -- main_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000001");
        state_var_NS <= main_C_1;
    END CASE;
  END PROCESS des_check_core_core_fsm_1;

  des_check_core_core_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= main_C_0;
      ELSE
        state_var <= state_var_NS;
      END IF;
    END IF;
  END PROCESS des_check_core_core_fsm_1_REG;

END v1;

-- ------------------------------------------------------------------
--  Design Unit:    des_check_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;


ENTITY des_check_core IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    input_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    input_rsc_triosy_lz : OUT STD_LOGIC;
    key_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    key_rsc_triosy_lz : OUT STD_LOGIC;
    return_rsc_dat : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    return_rsc_triosy_lz : OUT STD_LOGIC
  );
END des_check_core;

ARCHITECTURE v1 OF des_check_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL input_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL key_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL return_rsc_triosy_obj_ld : STD_LOGIC;
  SIGNAL return_rsci_idat_63 : STD_LOGIC;
  SIGNAL return_rsci_idat_62 : STD_LOGIC;
  SIGNAL return_rsci_idat_61 : STD_LOGIC;
  SIGNAL return_rsci_idat_60 : STD_LOGIC;
  SIGNAL return_rsci_idat_59 : STD_LOGIC;
  SIGNAL return_rsci_idat_58 : STD_LOGIC;
  SIGNAL return_rsci_idat_57 : STD_LOGIC;
  SIGNAL return_rsci_idat_56 : STD_LOGIC;
  SIGNAL return_rsci_idat_55 : STD_LOGIC;
  SIGNAL return_rsci_idat_54 : STD_LOGIC;
  SIGNAL return_rsci_idat_53 : STD_LOGIC;
  SIGNAL return_rsci_idat_52 : STD_LOGIC;
  SIGNAL return_rsci_idat_51 : STD_LOGIC;
  SIGNAL return_rsci_idat_50 : STD_LOGIC;
  SIGNAL return_rsci_idat_49 : STD_LOGIC;
  SIGNAL return_rsci_idat_48 : STD_LOGIC;
  SIGNAL return_rsci_idat_47 : STD_LOGIC;
  SIGNAL return_rsci_idat_46 : STD_LOGIC;
  SIGNAL return_rsci_idat_45 : STD_LOGIC;
  SIGNAL return_rsci_idat_44 : STD_LOGIC;
  SIGNAL return_rsci_idat_43 : STD_LOGIC;
  SIGNAL return_rsci_idat_42 : STD_LOGIC;
  SIGNAL return_rsci_idat_41 : STD_LOGIC;
  SIGNAL return_rsci_idat_40 : STD_LOGIC;
  SIGNAL return_rsci_idat_39 : STD_LOGIC;
  SIGNAL return_rsci_idat_38 : STD_LOGIC;
  SIGNAL return_rsci_idat_37 : STD_LOGIC;
  SIGNAL return_rsci_idat_36 : STD_LOGIC;
  SIGNAL return_rsci_idat_35 : STD_LOGIC;
  SIGNAL return_rsci_idat_34 : STD_LOGIC;
  SIGNAL return_rsci_idat_33 : STD_LOGIC;
  SIGNAL return_rsci_idat_32 : STD_LOGIC;
  SIGNAL return_rsci_idat_31 : STD_LOGIC;
  SIGNAL return_rsci_idat_30 : STD_LOGIC;
  SIGNAL return_rsci_idat_29 : STD_LOGIC;
  SIGNAL return_rsci_idat_28 : STD_LOGIC;
  SIGNAL return_rsci_idat_27 : STD_LOGIC;
  SIGNAL return_rsci_idat_26 : STD_LOGIC;
  SIGNAL return_rsci_idat_25 : STD_LOGIC;
  SIGNAL return_rsci_idat_24 : STD_LOGIC;
  SIGNAL return_rsci_idat_23 : STD_LOGIC;
  SIGNAL return_rsci_idat_22 : STD_LOGIC;
  SIGNAL return_rsci_idat_21 : STD_LOGIC;
  SIGNAL return_rsci_idat_20 : STD_LOGIC;
  SIGNAL return_rsci_idat_19 : STD_LOGIC;
  SIGNAL return_rsci_idat_18 : STD_LOGIC;
  SIGNAL return_rsci_idat_17 : STD_LOGIC;
  SIGNAL return_rsci_idat_16 : STD_LOGIC;
  SIGNAL return_rsci_idat_15 : STD_LOGIC;
  SIGNAL return_rsci_idat_14 : STD_LOGIC;
  SIGNAL return_rsci_idat_13 : STD_LOGIC;
  SIGNAL return_rsci_idat_12 : STD_LOGIC;
  SIGNAL return_rsci_idat_11 : STD_LOGIC;
  SIGNAL return_rsci_idat_10 : STD_LOGIC;
  SIGNAL return_rsci_idat_9 : STD_LOGIC;
  SIGNAL return_rsci_idat_8 : STD_LOGIC;
  SIGNAL return_rsci_idat_7 : STD_LOGIC;
  SIGNAL return_rsci_idat_6 : STD_LOGIC;
  SIGNAL return_rsci_idat_5 : STD_LOGIC;
  SIGNAL return_rsci_idat_4 : STD_LOGIC;
  SIGNAL return_rsci_idat_3 : STD_LOGIC;
  SIGNAL return_rsci_idat_2 : STD_LOGIC;
  SIGNAL return_rsci_idat_1 : STD_LOGIC;
  SIGNAL return_rsci_idat_0 : STD_LOGIC;
  SIGNAL fsm_output : STD_LOGIC_VECTOR (16 DOWNTO 0);
  SIGNAL reg_input_rsc_triosy_obj_ld_cse : STD_LOGIC;
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_6_itm : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_5_itm : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_2_itm : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_itm : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_1_itm : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_4_itm : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_3_itm : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_7_itm : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_14_itm : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_13_itm : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_10_itm : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_8_itm : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_9_itm : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_12_itm : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_11_itm : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_15_itm : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL input_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL key_io_read_key_rsc_cse_63_1_sva : STD_LOGIC_VECTOR (62 DOWNTO 0);
  SIGNAL s_output_1_19_16_19_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_23_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_34_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_38_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_49_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_53_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_4_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_8_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL R_15_1_sva : STD_LOGIC;
  SIGNAL R_16_1_sva : STD_LOGIC;
  SIGNAL R_14_1_sva : STD_LOGIC;
  SIGNAL R_17_1_sva : STD_LOGIC;
  SIGNAL R_13_1_sva : STD_LOGIC;
  SIGNAL R_18_1_sva : STD_LOGIC;
  SIGNAL R_12_1_sva : STD_LOGIC;
  SIGNAL R_19_1_sva : STD_LOGIC;
  SIGNAL R_11_1_sva : STD_LOGIC;
  SIGNAL R_20_1_sva : STD_LOGIC;
  SIGNAL R_10_1_sva : STD_LOGIC;
  SIGNAL R_21_1_sva : STD_LOGIC;
  SIGNAL R_9_1_sva : STD_LOGIC;
  SIGNAL R_22_1_sva : STD_LOGIC;
  SIGNAL R_8_1_sva : STD_LOGIC;
  SIGNAL R_23_1_sva : STD_LOGIC;
  SIGNAL R_7_1_sva : STD_LOGIC;
  SIGNAL R_24_1_sva : STD_LOGIC;
  SIGNAL R_6_1_sva : STD_LOGIC;
  SIGNAL R_25_1_sva : STD_LOGIC;
  SIGNAL R_5_1_sva : STD_LOGIC;
  SIGNAL R_26_1_sva : STD_LOGIC;
  SIGNAL R_4_1_sva : STD_LOGIC;
  SIGNAL R_27_1_sva : STD_LOGIC;
  SIGNAL R_3_1_sva : STD_LOGIC;
  SIGNAL R_28_1_sva : STD_LOGIC;
  SIGNAL R_2_1_sva : STD_LOGIC;
  SIGNAL R_29_1_sva : STD_LOGIC;
  SIGNAL R_1_1_sva : STD_LOGIC;
  SIGNAL R_30_1_sva : STD_LOGIC;
  SIGNAL R_0_1_sva : STD_LOGIC;
  SIGNAL R_31_1_sva : STD_LOGIC;
  SIGNAL s_output_1_19_16_20_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_24_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_35_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_39_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_50_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_54_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_5_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_9_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL R_15_3_sva : STD_LOGIC;
  SIGNAL R_16_3_sva : STD_LOGIC;
  SIGNAL R_14_3_sva : STD_LOGIC;
  SIGNAL R_17_3_sva : STD_LOGIC;
  SIGNAL R_13_3_sva : STD_LOGIC;
  SIGNAL R_18_3_sva : STD_LOGIC;
  SIGNAL R_12_3_sva : STD_LOGIC;
  SIGNAL R_19_3_sva : STD_LOGIC;
  SIGNAL R_11_3_sva : STD_LOGIC;
  SIGNAL R_20_3_sva : STD_LOGIC;
  SIGNAL R_10_3_sva : STD_LOGIC;
  SIGNAL R_21_3_sva : STD_LOGIC;
  SIGNAL R_9_3_sva : STD_LOGIC;
  SIGNAL R_22_3_sva : STD_LOGIC;
  SIGNAL R_8_3_sva : STD_LOGIC;
  SIGNAL R_23_3_sva : STD_LOGIC;
  SIGNAL R_7_3_sva : STD_LOGIC;
  SIGNAL R_24_3_sva : STD_LOGIC;
  SIGNAL R_6_3_sva : STD_LOGIC;
  SIGNAL R_25_3_sva : STD_LOGIC;
  SIGNAL R_5_3_sva : STD_LOGIC;
  SIGNAL R_26_3_sva : STD_LOGIC;
  SIGNAL R_4_3_sva : STD_LOGIC;
  SIGNAL R_27_3_sva : STD_LOGIC;
  SIGNAL R_3_3_sva : STD_LOGIC;
  SIGNAL R_28_3_sva : STD_LOGIC;
  SIGNAL R_2_3_sva : STD_LOGIC;
  SIGNAL R_29_3_sva : STD_LOGIC;
  SIGNAL R_1_3_sva : STD_LOGIC;
  SIGNAL R_30_3_sva : STD_LOGIC;
  SIGNAL R_0_3_sva : STD_LOGIC;
  SIGNAL R_31_3_sva : STD_LOGIC;
  SIGNAL R_15_4_sva : STD_LOGIC;
  SIGNAL R_16_4_sva : STD_LOGIC;
  SIGNAL R_14_4_sva : STD_LOGIC;
  SIGNAL R_17_4_sva : STD_LOGIC;
  SIGNAL R_13_4_sva : STD_LOGIC;
  SIGNAL R_18_4_sva : STD_LOGIC;
  SIGNAL R_12_4_sva : STD_LOGIC;
  SIGNAL R_19_4_sva : STD_LOGIC;
  SIGNAL R_11_4_sva : STD_LOGIC;
  SIGNAL R_20_4_sva : STD_LOGIC;
  SIGNAL R_10_4_sva : STD_LOGIC;
  SIGNAL R_21_4_sva : STD_LOGIC;
  SIGNAL R_9_4_sva : STD_LOGIC;
  SIGNAL R_22_4_sva : STD_LOGIC;
  SIGNAL R_8_4_sva : STD_LOGIC;
  SIGNAL R_23_4_sva : STD_LOGIC;
  SIGNAL R_7_4_sva : STD_LOGIC;
  SIGNAL R_24_4_sva : STD_LOGIC;
  SIGNAL R_6_4_sva : STD_LOGIC;
  SIGNAL R_25_4_sva : STD_LOGIC;
  SIGNAL R_5_4_sva : STD_LOGIC;
  SIGNAL R_26_4_sva : STD_LOGIC;
  SIGNAL R_4_4_sva : STD_LOGIC;
  SIGNAL R_27_4_sva : STD_LOGIC;
  SIGNAL R_3_4_sva : STD_LOGIC;
  SIGNAL R_28_4_sva : STD_LOGIC;
  SIGNAL R_2_4_sva : STD_LOGIC;
  SIGNAL R_29_4_sva : STD_LOGIC;
  SIGNAL R_1_4_sva : STD_LOGIC;
  SIGNAL R_30_4_sva : STD_LOGIC;
  SIGNAL R_0_4_sva : STD_LOGIC;
  SIGNAL R_31_4_sva : STD_LOGIC;
  SIGNAL R_15_5_sva : STD_LOGIC;
  SIGNAL R_16_5_sva : STD_LOGIC;
  SIGNAL R_14_5_sva : STD_LOGIC;
  SIGNAL R_17_5_sva : STD_LOGIC;
  SIGNAL R_13_5_sva : STD_LOGIC;
  SIGNAL R_18_5_sva : STD_LOGIC;
  SIGNAL R_12_5_sva : STD_LOGIC;
  SIGNAL R_19_5_sva : STD_LOGIC;
  SIGNAL R_11_5_sva : STD_LOGIC;
  SIGNAL R_20_5_sva : STD_LOGIC;
  SIGNAL R_10_5_sva : STD_LOGIC;
  SIGNAL R_21_5_sva : STD_LOGIC;
  SIGNAL R_9_5_sva : STD_LOGIC;
  SIGNAL R_22_5_sva : STD_LOGIC;
  SIGNAL R_8_5_sva : STD_LOGIC;
  SIGNAL R_23_5_sva : STD_LOGIC;
  SIGNAL R_7_5_sva : STD_LOGIC;
  SIGNAL R_24_5_sva : STD_LOGIC;
  SIGNAL R_6_5_sva : STD_LOGIC;
  SIGNAL R_25_5_sva : STD_LOGIC;
  SIGNAL R_5_5_sva : STD_LOGIC;
  SIGNAL R_26_5_sva : STD_LOGIC;
  SIGNAL R_4_5_sva : STD_LOGIC;
  SIGNAL R_27_5_sva : STD_LOGIC;
  SIGNAL R_3_5_sva : STD_LOGIC;
  SIGNAL R_28_5_sva : STD_LOGIC;
  SIGNAL R_2_5_sva : STD_LOGIC;
  SIGNAL R_29_5_sva : STD_LOGIC;
  SIGNAL R_1_5_sva : STD_LOGIC;
  SIGNAL R_30_5_sva : STD_LOGIC;
  SIGNAL R_0_5_sva : STD_LOGIC;
  SIGNAL R_31_5_sva : STD_LOGIC;
  SIGNAL R_15_6_sva : STD_LOGIC;
  SIGNAL R_16_6_sva : STD_LOGIC;
  SIGNAL R_14_6_sva : STD_LOGIC;
  SIGNAL R_17_6_sva : STD_LOGIC;
  SIGNAL R_13_6_sva : STD_LOGIC;
  SIGNAL R_18_6_sva : STD_LOGIC;
  SIGNAL R_12_6_sva : STD_LOGIC;
  SIGNAL R_19_6_sva : STD_LOGIC;
  SIGNAL R_11_6_sva : STD_LOGIC;
  SIGNAL R_20_6_sva : STD_LOGIC;
  SIGNAL R_10_6_sva : STD_LOGIC;
  SIGNAL R_21_6_sva : STD_LOGIC;
  SIGNAL R_9_6_sva : STD_LOGIC;
  SIGNAL R_22_6_sva : STD_LOGIC;
  SIGNAL R_8_6_sva : STD_LOGIC;
  SIGNAL R_23_6_sva : STD_LOGIC;
  SIGNAL R_7_6_sva : STD_LOGIC;
  SIGNAL R_24_6_sva : STD_LOGIC;
  SIGNAL R_6_6_sva : STD_LOGIC;
  SIGNAL R_25_6_sva : STD_LOGIC;
  SIGNAL R_5_6_sva : STD_LOGIC;
  SIGNAL R_26_6_sva : STD_LOGIC;
  SIGNAL R_4_6_sva : STD_LOGIC;
  SIGNAL R_27_6_sva : STD_LOGIC;
  SIGNAL R_3_6_sva : STD_LOGIC;
  SIGNAL R_28_6_sva : STD_LOGIC;
  SIGNAL R_2_6_sva : STD_LOGIC;
  SIGNAL R_29_6_sva : STD_LOGIC;
  SIGNAL R_1_6_sva : STD_LOGIC;
  SIGNAL R_30_6_sva : STD_LOGIC;
  SIGNAL R_0_6_sva : STD_LOGIC;
  SIGNAL R_31_6_sva : STD_LOGIC;
  SIGNAL R_15_7_sva : STD_LOGIC;
  SIGNAL R_16_7_sva : STD_LOGIC;
  SIGNAL R_14_7_sva : STD_LOGIC;
  SIGNAL R_17_7_sva : STD_LOGIC;
  SIGNAL R_13_7_sva : STD_LOGIC;
  SIGNAL R_18_7_sva : STD_LOGIC;
  SIGNAL R_12_7_sva : STD_LOGIC;
  SIGNAL R_19_7_sva : STD_LOGIC;
  SIGNAL R_11_7_sva : STD_LOGIC;
  SIGNAL R_20_7_sva : STD_LOGIC;
  SIGNAL R_10_7_sva : STD_LOGIC;
  SIGNAL R_21_7_sva : STD_LOGIC;
  SIGNAL R_9_7_sva : STD_LOGIC;
  SIGNAL R_22_7_sva : STD_LOGIC;
  SIGNAL R_8_7_sva : STD_LOGIC;
  SIGNAL R_23_7_sva : STD_LOGIC;
  SIGNAL R_7_7_sva : STD_LOGIC;
  SIGNAL R_24_7_sva : STD_LOGIC;
  SIGNAL R_6_7_sva : STD_LOGIC;
  SIGNAL R_25_7_sva : STD_LOGIC;
  SIGNAL R_5_7_sva : STD_LOGIC;
  SIGNAL R_26_7_sva : STD_LOGIC;
  SIGNAL R_4_7_sva : STD_LOGIC;
  SIGNAL R_27_7_sva : STD_LOGIC;
  SIGNAL R_3_7_sva : STD_LOGIC;
  SIGNAL R_28_7_sva : STD_LOGIC;
  SIGNAL R_2_7_sva : STD_LOGIC;
  SIGNAL R_29_7_sva : STD_LOGIC;
  SIGNAL R_1_7_sva : STD_LOGIC;
  SIGNAL R_30_7_sva : STD_LOGIC;
  SIGNAL R_0_7_sva : STD_LOGIC;
  SIGNAL R_31_7_sva : STD_LOGIC;
  SIGNAL R_15_8_sva : STD_LOGIC;
  SIGNAL R_16_8_sva : STD_LOGIC;
  SIGNAL R_14_8_sva : STD_LOGIC;
  SIGNAL R_17_8_sva : STD_LOGIC;
  SIGNAL R_13_8_sva : STD_LOGIC;
  SIGNAL R_18_8_sva : STD_LOGIC;
  SIGNAL R_12_8_sva : STD_LOGIC;
  SIGNAL R_19_8_sva : STD_LOGIC;
  SIGNAL R_11_8_sva : STD_LOGIC;
  SIGNAL R_20_8_sva : STD_LOGIC;
  SIGNAL R_10_8_sva : STD_LOGIC;
  SIGNAL R_21_8_sva : STD_LOGIC;
  SIGNAL R_9_8_sva : STD_LOGIC;
  SIGNAL R_22_8_sva : STD_LOGIC;
  SIGNAL R_8_8_sva : STD_LOGIC;
  SIGNAL R_23_8_sva : STD_LOGIC;
  SIGNAL R_7_8_sva : STD_LOGIC;
  SIGNAL R_24_8_sva : STD_LOGIC;
  SIGNAL R_6_8_sva : STD_LOGIC;
  SIGNAL R_25_8_sva : STD_LOGIC;
  SIGNAL R_5_8_sva : STD_LOGIC;
  SIGNAL R_26_8_sva : STD_LOGIC;
  SIGNAL R_4_8_sva : STD_LOGIC;
  SIGNAL R_27_8_sva : STD_LOGIC;
  SIGNAL R_3_8_sva : STD_LOGIC;
  SIGNAL R_28_8_sva : STD_LOGIC;
  SIGNAL R_2_8_sva : STD_LOGIC;
  SIGNAL R_29_8_sva : STD_LOGIC;
  SIGNAL R_1_8_sva : STD_LOGIC;
  SIGNAL R_30_8_sva : STD_LOGIC;
  SIGNAL R_0_8_sva : STD_LOGIC;
  SIGNAL R_31_8_sva : STD_LOGIC;
  SIGNAL R_15_9_sva : STD_LOGIC;
  SIGNAL R_16_9_sva : STD_LOGIC;
  SIGNAL R_14_9_sva : STD_LOGIC;
  SIGNAL R_17_9_sva : STD_LOGIC;
  SIGNAL R_13_9_sva : STD_LOGIC;
  SIGNAL R_18_9_sva : STD_LOGIC;
  SIGNAL R_12_9_sva : STD_LOGIC;
  SIGNAL R_19_9_sva : STD_LOGIC;
  SIGNAL R_11_9_sva : STD_LOGIC;
  SIGNAL R_20_9_sva : STD_LOGIC;
  SIGNAL R_10_9_sva : STD_LOGIC;
  SIGNAL R_21_9_sva : STD_LOGIC;
  SIGNAL R_9_9_sva : STD_LOGIC;
  SIGNAL R_22_9_sva : STD_LOGIC;
  SIGNAL R_8_9_sva : STD_LOGIC;
  SIGNAL R_23_9_sva : STD_LOGIC;
  SIGNAL R_7_9_sva : STD_LOGIC;
  SIGNAL R_24_9_sva : STD_LOGIC;
  SIGNAL R_6_9_sva : STD_LOGIC;
  SIGNAL R_25_9_sva : STD_LOGIC;
  SIGNAL R_5_9_sva : STD_LOGIC;
  SIGNAL R_26_9_sva : STD_LOGIC;
  SIGNAL R_4_9_sva : STD_LOGIC;
  SIGNAL R_27_9_sva : STD_LOGIC;
  SIGNAL R_3_9_sva : STD_LOGIC;
  SIGNAL R_28_9_sva : STD_LOGIC;
  SIGNAL R_2_9_sva : STD_LOGIC;
  SIGNAL R_29_9_sva : STD_LOGIC;
  SIGNAL R_1_9_sva : STD_LOGIC;
  SIGNAL R_30_9_sva : STD_LOGIC;
  SIGNAL R_0_9_sva : STD_LOGIC;
  SIGNAL R_31_9_sva : STD_LOGIC;
  SIGNAL R_15_10_sva : STD_LOGIC;
  SIGNAL R_16_10_sva : STD_LOGIC;
  SIGNAL R_14_10_sva : STD_LOGIC;
  SIGNAL R_17_10_sva : STD_LOGIC;
  SIGNAL R_13_10_sva : STD_LOGIC;
  SIGNAL R_18_10_sva : STD_LOGIC;
  SIGNAL R_12_10_sva : STD_LOGIC;
  SIGNAL R_19_10_sva : STD_LOGIC;
  SIGNAL R_11_10_sva : STD_LOGIC;
  SIGNAL R_20_10_sva : STD_LOGIC;
  SIGNAL R_10_10_sva : STD_LOGIC;
  SIGNAL R_21_10_sva : STD_LOGIC;
  SIGNAL R_9_10_sva : STD_LOGIC;
  SIGNAL R_22_10_sva : STD_LOGIC;
  SIGNAL R_8_10_sva : STD_LOGIC;
  SIGNAL R_23_10_sva : STD_LOGIC;
  SIGNAL R_7_10_sva : STD_LOGIC;
  SIGNAL R_24_10_sva : STD_LOGIC;
  SIGNAL R_6_10_sva : STD_LOGIC;
  SIGNAL R_25_10_sva : STD_LOGIC;
  SIGNAL R_5_10_sva : STD_LOGIC;
  SIGNAL R_26_10_sva : STD_LOGIC;
  SIGNAL R_4_10_sva : STD_LOGIC;
  SIGNAL R_27_10_sva : STD_LOGIC;
  SIGNAL R_3_10_sva : STD_LOGIC;
  SIGNAL R_28_10_sva : STD_LOGIC;
  SIGNAL R_2_10_sva : STD_LOGIC;
  SIGNAL R_29_10_sva : STD_LOGIC;
  SIGNAL R_1_10_sva : STD_LOGIC;
  SIGNAL R_30_10_sva : STD_LOGIC;
  SIGNAL R_0_10_sva : STD_LOGIC;
  SIGNAL R_31_10_sva : STD_LOGIC;
  SIGNAL R_15_11_sva : STD_LOGIC;
  SIGNAL R_16_11_sva : STD_LOGIC;
  SIGNAL R_14_11_sva : STD_LOGIC;
  SIGNAL R_17_11_sva : STD_LOGIC;
  SIGNAL R_13_11_sva : STD_LOGIC;
  SIGNAL R_18_11_sva : STD_LOGIC;
  SIGNAL R_12_11_sva : STD_LOGIC;
  SIGNAL R_19_11_sva : STD_LOGIC;
  SIGNAL R_11_11_sva : STD_LOGIC;
  SIGNAL R_20_11_sva : STD_LOGIC;
  SIGNAL R_10_11_sva : STD_LOGIC;
  SIGNAL R_21_11_sva : STD_LOGIC;
  SIGNAL R_9_11_sva : STD_LOGIC;
  SIGNAL R_22_11_sva : STD_LOGIC;
  SIGNAL R_8_11_sva : STD_LOGIC;
  SIGNAL R_23_11_sva : STD_LOGIC;
  SIGNAL R_7_11_sva : STD_LOGIC;
  SIGNAL R_24_11_sva : STD_LOGIC;
  SIGNAL R_6_11_sva : STD_LOGIC;
  SIGNAL R_25_11_sva : STD_LOGIC;
  SIGNAL R_5_11_sva : STD_LOGIC;
  SIGNAL R_26_11_sva : STD_LOGIC;
  SIGNAL R_4_11_sva : STD_LOGIC;
  SIGNAL R_27_11_sva : STD_LOGIC;
  SIGNAL R_3_11_sva : STD_LOGIC;
  SIGNAL R_28_11_sva : STD_LOGIC;
  SIGNAL R_2_11_sva : STD_LOGIC;
  SIGNAL R_29_11_sva : STD_LOGIC;
  SIGNAL R_1_11_sva : STD_LOGIC;
  SIGNAL R_30_11_sva : STD_LOGIC;
  SIGNAL R_0_11_sva : STD_LOGIC;
  SIGNAL R_31_11_sva : STD_LOGIC;
  SIGNAL R_15_12_sva : STD_LOGIC;
  SIGNAL R_16_12_sva : STD_LOGIC;
  SIGNAL R_14_12_sva : STD_LOGIC;
  SIGNAL R_17_12_sva : STD_LOGIC;
  SIGNAL R_13_12_sva : STD_LOGIC;
  SIGNAL R_18_12_sva : STD_LOGIC;
  SIGNAL R_12_12_sva : STD_LOGIC;
  SIGNAL R_19_12_sva : STD_LOGIC;
  SIGNAL R_11_12_sva : STD_LOGIC;
  SIGNAL R_20_12_sva : STD_LOGIC;
  SIGNAL R_10_12_sva : STD_LOGIC;
  SIGNAL R_21_12_sva : STD_LOGIC;
  SIGNAL R_9_12_sva : STD_LOGIC;
  SIGNAL R_22_12_sva : STD_LOGIC;
  SIGNAL R_8_12_sva : STD_LOGIC;
  SIGNAL R_23_12_sva : STD_LOGIC;
  SIGNAL R_7_12_sva : STD_LOGIC;
  SIGNAL R_24_12_sva : STD_LOGIC;
  SIGNAL R_6_12_sva : STD_LOGIC;
  SIGNAL R_25_12_sva : STD_LOGIC;
  SIGNAL R_5_12_sva : STD_LOGIC;
  SIGNAL R_26_12_sva : STD_LOGIC;
  SIGNAL R_4_12_sva : STD_LOGIC;
  SIGNAL R_27_12_sva : STD_LOGIC;
  SIGNAL R_3_12_sva : STD_LOGIC;
  SIGNAL R_28_12_sva : STD_LOGIC;
  SIGNAL R_2_12_sva : STD_LOGIC;
  SIGNAL R_29_12_sva : STD_LOGIC;
  SIGNAL R_1_12_sva : STD_LOGIC;
  SIGNAL R_30_12_sva : STD_LOGIC;
  SIGNAL R_0_12_sva : STD_LOGIC;
  SIGNAL R_31_12_sva : STD_LOGIC;
  SIGNAL R_15_13_sva : STD_LOGIC;
  SIGNAL R_16_13_sva : STD_LOGIC;
  SIGNAL R_14_13_sva : STD_LOGIC;
  SIGNAL R_17_13_sva : STD_LOGIC;
  SIGNAL R_13_13_sva : STD_LOGIC;
  SIGNAL R_18_13_sva : STD_LOGIC;
  SIGNAL R_12_13_sva : STD_LOGIC;
  SIGNAL R_19_13_sva : STD_LOGIC;
  SIGNAL R_11_13_sva : STD_LOGIC;
  SIGNAL R_20_13_sva : STD_LOGIC;
  SIGNAL R_10_13_sva : STD_LOGIC;
  SIGNAL R_21_13_sva : STD_LOGIC;
  SIGNAL R_9_13_sva : STD_LOGIC;
  SIGNAL R_22_13_sva : STD_LOGIC;
  SIGNAL R_8_13_sva : STD_LOGIC;
  SIGNAL R_23_13_sva : STD_LOGIC;
  SIGNAL R_7_13_sva : STD_LOGIC;
  SIGNAL R_24_13_sva : STD_LOGIC;
  SIGNAL R_6_13_sva : STD_LOGIC;
  SIGNAL R_25_13_sva : STD_LOGIC;
  SIGNAL R_5_13_sva : STD_LOGIC;
  SIGNAL R_26_13_sva : STD_LOGIC;
  SIGNAL R_4_13_sva : STD_LOGIC;
  SIGNAL R_27_13_sva : STD_LOGIC;
  SIGNAL R_3_13_sva : STD_LOGIC;
  SIGNAL R_28_13_sva : STD_LOGIC;
  SIGNAL R_2_13_sva : STD_LOGIC;
  SIGNAL R_29_13_sva : STD_LOGIC;
  SIGNAL R_1_13_sva : STD_LOGIC;
  SIGNAL R_30_13_sva : STD_LOGIC;
  SIGNAL R_0_13_sva : STD_LOGIC;
  SIGNAL R_31_13_sva : STD_LOGIC;
  SIGNAL R_15_14_sva : STD_LOGIC;
  SIGNAL R_16_14_sva : STD_LOGIC;
  SIGNAL R_14_14_sva : STD_LOGIC;
  SIGNAL R_17_14_sva : STD_LOGIC;
  SIGNAL R_13_14_sva : STD_LOGIC;
  SIGNAL R_18_14_sva : STD_LOGIC;
  SIGNAL R_12_14_sva : STD_LOGIC;
  SIGNAL R_19_14_sva : STD_LOGIC;
  SIGNAL R_11_14_sva : STD_LOGIC;
  SIGNAL R_20_14_sva : STD_LOGIC;
  SIGNAL R_10_14_sva : STD_LOGIC;
  SIGNAL R_21_14_sva : STD_LOGIC;
  SIGNAL R_9_14_sva : STD_LOGIC;
  SIGNAL R_22_14_sva : STD_LOGIC;
  SIGNAL R_8_14_sva : STD_LOGIC;
  SIGNAL R_23_14_sva : STD_LOGIC;
  SIGNAL R_7_14_sva : STD_LOGIC;
  SIGNAL R_24_14_sva : STD_LOGIC;
  SIGNAL R_6_14_sva : STD_LOGIC;
  SIGNAL R_25_14_sva : STD_LOGIC;
  SIGNAL R_5_14_sva : STD_LOGIC;
  SIGNAL R_26_14_sva : STD_LOGIC;
  SIGNAL R_4_14_sva : STD_LOGIC;
  SIGNAL R_27_14_sva : STD_LOGIC;
  SIGNAL R_3_14_sva : STD_LOGIC;
  SIGNAL R_28_14_sva : STD_LOGIC;
  SIGNAL R_2_14_sva : STD_LOGIC;
  SIGNAL R_29_14_sva : STD_LOGIC;
  SIGNAL R_1_14_sva : STD_LOGIC;
  SIGNAL R_30_14_sva : STD_LOGIC;
  SIGNAL R_0_14_sva : STD_LOGIC;
  SIGNAL R_31_14_sva : STD_LOGIC;
  SIGNAL R_15_15_sva : STD_LOGIC;
  SIGNAL R_16_15_sva : STD_LOGIC;
  SIGNAL R_14_15_sva : STD_LOGIC;
  SIGNAL R_17_15_sva : STD_LOGIC;
  SIGNAL R_13_15_sva : STD_LOGIC;
  SIGNAL R_18_15_sva : STD_LOGIC;
  SIGNAL R_12_15_sva : STD_LOGIC;
  SIGNAL R_19_15_sva : STD_LOGIC;
  SIGNAL R_11_15_sva : STD_LOGIC;
  SIGNAL R_20_15_sva : STD_LOGIC;
  SIGNAL R_10_15_sva : STD_LOGIC;
  SIGNAL R_21_15_sva : STD_LOGIC;
  SIGNAL R_9_15_sva : STD_LOGIC;
  SIGNAL R_22_15_sva : STD_LOGIC;
  SIGNAL R_8_15_sva : STD_LOGIC;
  SIGNAL R_23_15_sva : STD_LOGIC;
  SIGNAL R_7_15_sva : STD_LOGIC;
  SIGNAL R_24_15_sva : STD_LOGIC;
  SIGNAL R_6_15_sva : STD_LOGIC;
  SIGNAL R_25_15_sva : STD_LOGIC;
  SIGNAL R_5_15_sva : STD_LOGIC;
  SIGNAL R_26_15_sva : STD_LOGIC;
  SIGNAL R_4_15_sva : STD_LOGIC;
  SIGNAL R_27_15_sva : STD_LOGIC;
  SIGNAL R_3_15_sva : STD_LOGIC;
  SIGNAL R_28_15_sva : STD_LOGIC;
  SIGNAL R_2_15_sva : STD_LOGIC;
  SIGNAL R_29_15_sva : STD_LOGIC;
  SIGNAL R_1_15_sva : STD_LOGIC;
  SIGNAL R_30_15_sva : STD_LOGIC;
  SIGNAL R_0_15_sva : STD_LOGIC;
  SIGNAL R_31_15_sva : STD_LOGIC;
  SIGNAL s_output_1_19_16_6_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_55_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_36_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_21_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_25_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_51_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_40_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_10_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_7_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_56_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_37_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_22_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_26_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_52_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_41_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_11_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_8_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_57_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_38_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_23_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_27_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_53_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_42_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_12_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_9_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_58_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_39_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_24_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_28_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_54_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_43_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_13_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_10_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_59_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_40_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_25_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_29_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_55_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_44_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_14_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_11_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_60_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_41_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_26_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_30_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_56_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_45_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_15_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_12_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_61_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_42_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_27_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_31_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_57_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_46_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_16_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_13_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_62_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_43_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_28_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_32_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_58_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_47_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_17_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_14_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_63_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_44_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_29_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_33_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_59_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_48_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_18_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_15_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_64_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_45_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_30_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_34_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_60_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_49_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_19_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_16_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_65_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_46_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_31_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_35_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_61_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_50_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_20_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_17_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_66_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_47_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_32_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_36_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_62_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_51_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_21_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_18_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_67_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_48_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_33_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_37_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_63_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_52_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_22_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_5_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_1_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_3_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_7_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_19_16_2_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL s_output_1_3_0_6_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL loop_DES_rounds_1_xor_32_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_32_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_31_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_31_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_30_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_30_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_29_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_29_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_28_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_28_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_27_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_27_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_26_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_26_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_25_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_25_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_24_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_24_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_23_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_23_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_22_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_22_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_21_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_21_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_20_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_20_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_19_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_19_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_18_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_18_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_17_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_17_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_16_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_16_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_15_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_15_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_14_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_14_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_13_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_13_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_12_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_12_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_11_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_11_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_10_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_10_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_9_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_9_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_8_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_8_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_7_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_7_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_6_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_6_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_5_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_5_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_4_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_4_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_3_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_3_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_2_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_2_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_1_xor_1_nl : STD_LOGIC;
  SIGNAL loop_DES_rounds_2_xor_1_nl : STD_LOGIC;
  SIGNAL input_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL input_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL key_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL key_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL return_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL return_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_6_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_6_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_5_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_5_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_2_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_2_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_rg_addr : STD_LOGIC_VECTOR (8 DOWNTO
      0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_rg_data_out : STD_LOGIC_VECTOR (3
      DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_1_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_1_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_4_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_4_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_3_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_3_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_7_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_7_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_14_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_14_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_13_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_13_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_10_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_10_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_8_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_8_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_9_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_9_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_12_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_12_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_11_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_11_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_15_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_15_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_22_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_22_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_21_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_21_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_18_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_18_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_16_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_16_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_17_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_17_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_20_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_20_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_19_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_19_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_23_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_23_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_30_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_30_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_29_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_29_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_26_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_26_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_24_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_24_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_25_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_25_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_28_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_28_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_27_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_27_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_31_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_31_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_38_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_38_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_37_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_37_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_34_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_34_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_32_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_32_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_33_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_33_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_36_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_36_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_35_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_35_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_39_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_39_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_46_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_46_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_45_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_45_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_42_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_42_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_40_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_40_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_41_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_41_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_44_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_44_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_43_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_43_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_47_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_47_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_54_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_54_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_53_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_53_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_50_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_50_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_48_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_48_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_49_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_49_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_52_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_52_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_51_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_51_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_55_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_55_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_62_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_62_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_61_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_61_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_58_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_58_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_56_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_56_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_57_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_57_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_60_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_60_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_59_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_59_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_63_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_63_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_70_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_70_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_69_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_69_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_66_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_66_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_64_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_64_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_65_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_65_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_68_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_68_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_67_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_67_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_71_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_71_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_78_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_78_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_77_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_77_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_74_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_74_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_72_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_72_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_73_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_73_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_76_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_76_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_75_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_75_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_79_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_79_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_86_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_86_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_85_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_85_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_82_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_82_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_80_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_80_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_81_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_81_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_84_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_84_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_83_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_83_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_87_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_87_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_94_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_94_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_93_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_93_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_90_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_90_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_88_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_88_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_89_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_89_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_92_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_92_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_91_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_91_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_95_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_95_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_102_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_102_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_101_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_101_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_98_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_98_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_96_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_96_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_97_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_97_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_100_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_100_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_99_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_99_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_103_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_103_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_110_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_110_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_109_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_109_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_106_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_106_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_104_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_104_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_105_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_105_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_108_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_108_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_107_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_107_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_111_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_111_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_118_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_118_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_117_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_117_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_114_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_114_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_112_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_112_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_113_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_113_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_116_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_116_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_115_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_115_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_119_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_119_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_121_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_121_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_120_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_120_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_124_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_124_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_126_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_126_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_125_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_125_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_122_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_122_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_127_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_127_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_123_rg_addr : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL operator_8_false_1_read_rom_S_rom_map_1_123_rg_data_out : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

  COMPONENT des_check_core_core_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (16 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL des_check_core_core_fsm_inst_fsm_output : STD_LOGIC_VECTOR (16 DOWNTO 0);

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  input_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 1,
      width => 64
      )
    PORT MAP(
      dat => input_rsci_dat,
      idat => input_rsci_idat_1
    );
  input_rsci_dat <= input_rsc_dat;
  input_rsci_idat <= input_rsci_idat_1;

  key_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 2,
      width => 64
      )
    PORT MAP(
      dat => key_rsci_dat,
      idat => key_rsci_idat_1
    );
  key_rsci_dat <= key_rsc_dat;
  key_rsci_idat <= key_rsci_idat_1;

  return_rsci : work.ccs_out_pkg_v1.ccs_out_v1
    GENERIC MAP(
      rscid => 3,
      width => 64
      )
    PORT MAP(
      idat => return_rsci_idat,
      dat => return_rsci_dat
    );
  return_rsci_idat <= STD_LOGIC_VECTOR'( return_rsci_idat_63 & return_rsci_idat_62
      & return_rsci_idat_61 & return_rsci_idat_60 & return_rsci_idat_59 & return_rsci_idat_58
      & return_rsci_idat_57 & return_rsci_idat_56 & return_rsci_idat_55 & return_rsci_idat_54
      & return_rsci_idat_53 & return_rsci_idat_52 & return_rsci_idat_51 & return_rsci_idat_50
      & return_rsci_idat_49 & return_rsci_idat_48 & return_rsci_idat_47 & return_rsci_idat_46
      & return_rsci_idat_45 & return_rsci_idat_44 & return_rsci_idat_43 & return_rsci_idat_42
      & return_rsci_idat_41 & return_rsci_idat_40 & return_rsci_idat_39 & return_rsci_idat_38
      & return_rsci_idat_37 & return_rsci_idat_36 & return_rsci_idat_35 & return_rsci_idat_34
      & return_rsci_idat_33 & return_rsci_idat_32 & return_rsci_idat_31 & return_rsci_idat_30
      & return_rsci_idat_29 & return_rsci_idat_28 & return_rsci_idat_27 & return_rsci_idat_26
      & return_rsci_idat_25 & return_rsci_idat_24 & return_rsci_idat_23 & return_rsci_idat_22
      & return_rsci_idat_21 & return_rsci_idat_20 & return_rsci_idat_19 & return_rsci_idat_18
      & return_rsci_idat_17 & return_rsci_idat_16 & return_rsci_idat_15 & return_rsci_idat_14
      & return_rsci_idat_13 & return_rsci_idat_12 & return_rsci_idat_11 & return_rsci_idat_10
      & return_rsci_idat_9 & return_rsci_idat_8 & return_rsci_idat_7 & return_rsci_idat_6
      & return_rsci_idat_5 & return_rsci_idat_4 & return_rsci_idat_3 & return_rsci_idat_2
      & return_rsci_idat_1 & return_rsci_idat_0);
  return_rsc_dat <= return_rsci_dat;

  input_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_input_rsc_triosy_obj_ld_cse,
      lz => input_rsc_triosy_lz
    );
  key_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_input_rsc_triosy_obj_ld_cse,
      lz => key_rsc_triosy_lz
    );
  return_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => return_rsc_triosy_obj_ld,
      lz => return_rsc_triosy_lz
    );
  operator_8_false_1_read_rom_S_rom_map_1_6_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_6_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_6_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_6_rg_addr <= STD_LOGIC_VECTOR'( "011")
      & ((input_rsci_idat(29)) XOR (key_rsci_idat(5))) & ((input_rsci_idat(3)) XOR
      (key_rsci_idat(23))) & ((input_rsci_idat(37)) XOR (key_rsci_idat(63))) & ((input_rsci_idat(45))
      XOR (key_rsci_idat(28))) & ((input_rsci_idat(53)) XOR (key_rsci_idat(37)))
      & ((input_rsci_idat(61)) XOR (key_rsci_idat(46)));
  operator_8_false_1_read_rom_S_rom_map_1_6_itm <= operator_8_false_1_read_rom_S_rom_map_1_6_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_5_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_5_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_5_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_5_rg_addr <= STD_LOGIC_VECTOR'( "110")
      & ((input_rsci_idat(59)) XOR (key_rsci_idat(3))) & ((input_rsci_idat(33)) XOR
      (key_rsci_idat(44))) & ((input_rsci_idat(1)) XOR (key_rsci_idat(43))) & ((input_rsci_idat(9))
      XOR (key_rsci_idat(26))) & ((input_rsci_idat(17)) XOR (key_rsci_idat(1))) &
      ((input_rsci_idat(25)) XOR (key_rsci_idat(49)));
  operator_8_false_1_read_rom_S_rom_map_1_5_itm <= operator_8_false_1_read_rom_S_rom_map_1_5_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_2_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_2_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_2_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_2_rg_addr <= STD_LOGIC_VECTOR'( "001")
      & ((input_rsci_idat(31)) XOR (key_rsci_idat(31))) & ((input_rsci_idat(5)) XOR
      (key_rsci_idat(22))) & ((input_rsci_idat(39)) XOR (key_rsci_idat(7))) & ((input_rsci_idat(47))
      XOR (key_rsci_idat(62))) & ((input_rsci_idat(55)) XOR (key_rsci_idat(55)))
      & ((input_rsci_idat(63)) XOR (key_rsci_idat(45)));
  operator_8_false_1_read_rom_S_rom_map_1_2_itm <= operator_8_false_1_read_rom_S_rom_map_1_2_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_rg_addr <= STD_LOGIC_VECTOR'( "000") &
      ((input_rsci_idat(57)) XOR (key_rsci_idat(54))) & ((input_rsci_idat(39)) XOR
      (key_rsci_idat(47))) & ((input_rsci_idat(7)) XOR (key_rsci_idat(13))) & ((input_rsci_idat(15))
      XOR (key_rsci_idat(30))) & ((input_rsci_idat(23)) XOR (key_rsci_idat(4))) &
      ((input_rsci_idat(31)) XOR (key_rsci_idat(15)));
  operator_8_false_1_read_rom_S_rom_map_1_itm <= operator_8_false_1_read_rom_S_rom_map_1_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_1_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_1_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_1_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_1_rg_addr <= STD_LOGIC_VECTOR'( "100")
      & ((input_rsci_idat(61)) XOR (key_rsci_idat(42))) & ((input_rsci_idat(35))
      XOR (key_rsci_idat(60))) & ((input_rsci_idat(3)) XOR (key_rsci_idat(36))) &
      ((input_rsci_idat(11)) XOR (key_rsci_idat(25))) & ((input_rsci_idat(19)) XOR
      (key_rsci_idat(10))) & ((input_rsci_idat(27)) XOR (key_rsci_idat(27)));
  operator_8_false_1_read_rom_S_rom_map_1_1_itm <= operator_8_false_1_read_rom_S_rom_map_1_1_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_4_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_4_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_4_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_4_rg_addr <= STD_LOGIC_VECTOR'( "010")
      & ((input_rsci_idat(63)) XOR (key_rsci_idat(61))) & ((input_rsci_idat(37))
      XOR (key_rsci_idat(6))) & ((input_rsci_idat(5)) XOR (key_rsci_idat(29))) &
      ((input_rsci_idat(13)) XOR (key_rsci_idat(38))) & ((input_rsci_idat(21)) XOR
      (key_rsci_idat(39))) & ((input_rsci_idat(29)) XOR (key_rsci_idat(20)));
  operator_8_false_1_read_rom_S_rom_map_1_4_itm <= operator_8_false_1_read_rom_S_rom_map_1_4_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_3_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_3_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_3_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_3_rg_addr <= STD_LOGIC_VECTOR'( "101")
      & ((input_rsci_idat(27)) XOR (key_rsci_idat(17))) & ((input_rsci_idat(1)) XOR
      (key_rsci_idat(35))) & ((input_rsci_idat(35)) XOR (key_rsci_idat(34))) & ((input_rsci_idat(43))
      XOR (key_rsci_idat(59))) & ((input_rsci_idat(51)) XOR (key_rsci_idat(11)))
      & ((input_rsci_idat(59)) XOR (key_rsci_idat(41)));
  operator_8_false_1_read_rom_S_rom_map_1_3_itm <= operator_8_false_1_read_rom_S_rom_map_1_3_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_7_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_7_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_7_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_7_rg_addr <= STD_LOGIC_VECTOR'( "111")
      & ((input_rsci_idat(25)) XOR (key_rsci_idat(19))) & ((input_rsci_idat(7)) XOR
      (key_rsci_idat(33))) & ((input_rsci_idat(33)) XOR (key_rsci_idat(50))) & ((input_rsci_idat(41))
      XOR (key_rsci_idat(51))) & ((input_rsci_idat(49)) XOR (key_rsci_idat(2))) &
      ((input_rsci_idat(57)) XOR (key_rsci_idat(9)));
  operator_8_false_1_read_rom_S_rom_map_1_7_itm <= operator_8_false_1_read_rom_S_rom_map_1_7_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_14_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_14_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_14_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_14_rg_addr <= STD_LOGIC_VECTOR'( "011")
      & ((input_sva(28)) XOR (s_output_1_3_0_53_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(12)))
      & ((input_sva(2)) XOR (s_output_1_19_16_19_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(30)))
      & ((input_sva(36)) XOR (s_output_1_19_16_34_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(5)))
      & ((input_sva(44)) XOR (s_output_1_3_0_23_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(6)))
      & ((input_sva(52)) XOR (s_output_1_3_0_8_sva(1)) XOR (key_io_read_key_rsc_cse_63_1_sva(44)))
      & ((input_sva(60)) XOR (s_output_1_19_16_49_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(53)));
  operator_8_false_1_read_rom_S_rom_map_1_14_itm <= operator_8_false_1_read_rom_S_rom_map_1_14_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_13_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_13_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_13_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_13_rg_addr <= STD_LOGIC_VECTOR'( "110")
      & ((input_sva(58)) XOR (s_output_1_19_16_49_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(10)))
      & ((input_sva(32)) XOR (s_output_1_3_0_38_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(51)))
      & ((input_sva(0)) XOR (s_output_1_3_0_23_sva(1)) XOR (key_io_read_key_rsc_cse_63_1_sva(50)))
      & ((input_sva(8)) XOR (s_output_1_19_16_4_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(33)))
      & ((input_sva(16)) XOR (s_output_1_3_0_8_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(8)))
      & ((input_sva(24)) XOR (s_output_1_19_16_34_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(56)));
  operator_8_false_1_read_rom_S_rom_map_1_13_itm <= operator_8_false_1_read_rom_S_rom_map_1_13_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_10_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_10_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_10_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_10_rg_addr <= STD_LOGIC_VECTOR'( "001")
      & ((input_sva(30)) XOR (s_output_1_3_0_38_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(38)))
      & ((input_sva(4)) XOR (s_output_1_19_16_19_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(29)))
      & ((input_sva(38)) XOR (s_output_1_3_0_8_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(14)))
      & ((input_sva(46)) XOR (s_output_1_19_16_49_sva(0)) XOR (key_io_read_key_rsc_cse_63_1_sva(4)))
      & ((input_sva(54)) XOR (s_output_1_3_0_53_sva(0)) XOR (key_io_read_key_rsc_cse_63_1_sva(62)))
      & ((input_sva(62)) XOR (s_output_1_3_0_23_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(52)));
  operator_8_false_1_read_rom_S_rom_map_1_10_itm <= operator_8_false_1_read_rom_S_rom_map_1_10_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_8_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_8_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_8_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_8_rg_addr <= STD_LOGIC_VECTOR'( "000")
      & ((input_sva(56)) XOR (s_output_1_3_0_53_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(61)))
      & ((input_sva(38)) XOR (s_output_1_3_0_8_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(54)))
      & ((input_sva(6)) XOR (s_output_1_19_16_4_sva(0)) XOR (key_io_read_key_rsc_cse_63_1_sva(20)))
      & ((input_sva(14)) XOR (s_output_1_19_16_34_sva(1)) XOR (key_io_read_key_rsc_cse_63_1_sva(37)))
      & ((input_sva(22)) XOR (s_output_1_3_0_23_sva(0)) XOR (key_io_read_key_rsc_cse_63_1_sva(11)))
      & ((input_sva(30)) XOR (s_output_1_3_0_38_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(22)));
  operator_8_false_1_read_rom_S_rom_map_1_8_itm <= operator_8_false_1_read_rom_S_rom_map_1_8_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_9_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_9_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_9_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_9_rg_addr <= STD_LOGIC_VECTOR'( "100")
      & ((input_sva(60)) XOR (s_output_1_19_16_49_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(49)))
      & ((input_sva(34)) XOR (s_output_1_3_0_8_sva(0)) XOR (key_io_read_key_rsc_cse_63_1_sva(0)))
      & ((input_sva(2)) XOR (s_output_1_19_16_19_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(43)))
      & ((input_sva(10)) XOR (s_output_1_19_16_34_sva(0)) XOR (key_io_read_key_rsc_cse_63_1_sva(32)))
      & ((input_sva(18)) XOR (s_output_1_3_0_38_sva(0)) XOR (key_io_read_key_rsc_cse_63_1_sva(17)))
      & ((input_sva(26)) XOR (s_output_1_19_16_4_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(34)));
  operator_8_false_1_read_rom_S_rom_map_1_9_itm <= operator_8_false_1_read_rom_S_rom_map_1_9_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_12_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_12_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_12_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_12_rg_addr <= STD_LOGIC_VECTOR'( "010")
      & ((input_sva(62)) XOR (s_output_1_3_0_23_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(3)))
      & ((input_sva(36)) XOR (s_output_1_19_16_34_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(13)))
      & ((input_sva(4)) XOR (s_output_1_19_16_19_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(36)))
      & ((input_sva(12)) XOR (s_output_1_19_16_4_sva(1)) XOR (key_io_read_key_rsc_cse_63_1_sva(45)))
      & ((input_sva(20)) XOR (s_output_1_3_0_38_sva(1)) XOR (key_io_read_key_rsc_cse_63_1_sva(46)))
      & ((input_sva(28)) XOR (s_output_1_3_0_53_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(27)));
  operator_8_false_1_read_rom_S_rom_map_1_12_itm <= operator_8_false_1_read_rom_S_rom_map_1_12_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_11_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_11_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_11_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_11_rg_addr <= STD_LOGIC_VECTOR'( "101")
      & ((input_sva(26)) XOR (s_output_1_19_16_4_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(24)))
      & ((input_sva(0)) XOR (s_output_1_3_0_23_sva(1)) XOR (key_io_read_key_rsc_cse_63_1_sva(42)))
      & ((key_io_read_key_rsc_cse_63_1_sva(41)) XOR (input_sva(34)) XOR (s_output_1_3_0_8_sva(0)))
      & ((input_sva(42)) XOR (s_output_1_3_0_53_sva(1)) XOR (key_io_read_key_rsc_cse_63_1_sva(35)))
      & ((input_sva(50)) XOR (s_output_1_19_16_19_sva(1)) XOR (key_io_read_key_rsc_cse_63_1_sva(18)))
      & ((input_sva(58)) XOR (s_output_1_19_16_49_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(48)));
  operator_8_false_1_read_rom_S_rom_map_1_11_itm <= operator_8_false_1_read_rom_S_rom_map_1_11_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_15_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_15_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_15_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_15_rg_addr <= STD_LOGIC_VECTOR'( "111")
      & ((input_sva(24)) XOR (s_output_1_19_16_34_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(26)))
      & ((input_sva(6)) XOR (s_output_1_19_16_4_sva(0)) XOR (key_io_read_key_rsc_cse_63_1_sva(40)))
      & ((input_sva(32)) XOR (s_output_1_3_0_38_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(57)))
      & ((input_sva(40)) XOR (s_output_1_19_16_49_sva(1)) XOR (key_io_read_key_rsc_cse_63_1_sva(58)))
      & ((input_sva(48)) XOR (s_output_1_19_16_19_sva(0)) XOR (key_io_read_key_rsc_cse_63_1_sva(9)))
      & ((input_sva(56)) XOR (s_output_1_3_0_53_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(16)));
  operator_8_false_1_read_rom_S_rom_map_1_15_itm <= operator_8_false_1_read_rom_S_rom_map_1_15_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_22_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_22_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_22_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_22_rg_addr <= STD_LOGIC_VECTOR'( "011")
      & ((key_io_read_key_rsc_cse_63_1_sva(28)) XOR (input_sva(29)) XOR (s_output_1_3_0_54_sva(2)))
      & ((input_sva(3)) XOR (s_output_1_19_16_20_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(46)))
      & ((key_io_read_key_rsc_cse_63_1_sva(21)) XOR (input_sva(37)) XOR (s_output_1_19_16_35_sva(3)))
      & ((input_sva(45)) XOR (s_output_1_3_0_24_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(22)))
      & ((input_sva(53)) XOR (s_output_1_3_0_9_sva(1)) XOR (key_io_read_key_rsc_cse_63_1_sva(60)))
      & ((input_sva(61)) XOR (s_output_1_19_16_50_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(4)));
  s_output_1_19_16_6_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_22_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_21_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_21_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_21_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_21_rg_addr <= STD_LOGIC_VECTOR'( "110")
      & ((input_sva(59)) XOR (s_output_1_19_16_50_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(26)))
      & ((input_sva(33)) XOR (s_output_1_3_0_39_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(0)))
      & ((input_sva(1)) XOR (s_output_1_3_0_24_sva(1)) XOR (key_io_read_key_rsc_cse_63_1_sva(35)))
      & ((input_sva(9)) XOR (s_output_1_19_16_5_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(49)))
      & ((input_sva(17)) XOR (s_output_1_3_0_9_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(24)))
      & ((input_sva(25)) XOR (s_output_1_19_16_35_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(9)));
  s_output_1_3_0_55_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_21_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_18_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_18_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_18_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_18_rg_addr <= STD_LOGIC_VECTOR'( "001")
      & ((input_sva(31)) XOR (s_output_1_3_0_39_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(54)))
      & ((input_sva(5)) XOR (s_output_1_19_16_20_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(45)))
      & ((input_sva(39)) XOR (s_output_1_3_0_9_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(30)))
      & ((input_sva(47)) XOR (s_output_1_19_16_50_sva(0)) XOR (key_io_read_key_rsc_cse_63_1_sva(20)))
      & ((input_sva(55)) XOR (s_output_1_3_0_54_sva(0)) XOR (key_io_read_key_rsc_cse_63_1_sva(13)))
      & ((input_sva(63)) XOR (s_output_1_3_0_24_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(3)));
  s_output_1_19_16_36_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_18_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_16_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_16_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_16_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_16_rg_addr <= STD_LOGIC_VECTOR'( "000")
      & ((input_sva(57)) XOR (s_output_1_3_0_54_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(12)))
      & ((input_sva(39)) XOR (s_output_1_3_0_9_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(5)))
      & ((input_sva(7)) XOR (s_output_1_19_16_5_sva(0)) XOR (key_io_read_key_rsc_cse_63_1_sva(36)))
      & ((input_sva(15)) XOR (s_output_1_19_16_35_sva(1)) XOR (key_io_read_key_rsc_cse_63_1_sva(53)))
      & ((input_sva(23)) XOR (s_output_1_3_0_24_sva(0)) XOR (key_io_read_key_rsc_cse_63_1_sva(27)))
      & ((input_sva(31)) XOR (s_output_1_3_0_39_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(38)));
  s_output_1_19_16_21_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_16_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_17_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_17_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_17_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_17_rg_addr <= STD_LOGIC_VECTOR'( "100")
      & ((key_io_read_key_rsc_cse_63_1_sva(2)) XOR (input_sva(61)) XOR (s_output_1_19_16_50_sva(2)))
      & ((input_sva(35)) XOR (s_output_1_3_0_9_sva(0)) XOR (key_io_read_key_rsc_cse_63_1_sva(16)))
      & ((key_io_read_key_rsc_cse_63_1_sva(59)) XOR (input_sva(3)) XOR (s_output_1_19_16_20_sva(2)))
      & ((input_sva(11)) XOR (s_output_1_19_16_35_sva(0)) XOR (key_io_read_key_rsc_cse_63_1_sva(48)))
      & ((input_sva(19)) XOR (s_output_1_3_0_39_sva(0)) XOR (key_io_read_key_rsc_cse_63_1_sva(33)))
      & ((input_sva(27)) XOR (s_output_1_19_16_5_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(50)));
  s_output_1_3_0_25_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_17_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_20_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_20_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_20_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_20_rg_addr <= STD_LOGIC_VECTOR'( "010")
      & ((key_io_read_key_rsc_cse_63_1_sva(19)) XOR (input_sva(63)) XOR (s_output_1_3_0_24_sva(3)))
      & ((input_sva(37)) XOR (s_output_1_19_16_35_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(29)))
      & ((input_sva(5)) XOR (s_output_1_19_16_20_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(52)))
      & ((input_sva(13)) XOR (s_output_1_19_16_5_sva(1)) XOR (key_io_read_key_rsc_cse_63_1_sva(61)))
      & ((input_sva(21)) XOR (s_output_1_3_0_39_sva(1)) XOR (key_io_read_key_rsc_cse_63_1_sva(62)))
      & ((input_sva(29)) XOR (s_output_1_3_0_54_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(14)));
  s_output_1_19_16_51_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_20_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_19_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_19_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_19_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_19_rg_addr <= STD_LOGIC_VECTOR'( "101")
      & ((input_sva(27)) XOR (s_output_1_19_16_5_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(40)))
      & ((input_sva(1)) XOR (s_output_1_3_0_24_sva(1)) XOR (key_io_read_key_rsc_cse_63_1_sva(58)))
      & ((input_sva(35)) XOR (s_output_1_3_0_9_sva(0)) XOR (key_io_read_key_rsc_cse_63_1_sva(57)))
      & ((input_sva(43)) XOR (s_output_1_3_0_54_sva(1)) XOR (key_io_read_key_rsc_cse_63_1_sva(51)))
      & ((input_sva(51)) XOR (s_output_1_19_16_20_sva(1)) XOR (key_io_read_key_rsc_cse_63_1_sva(34)))
      & ((key_io_read_key_rsc_cse_63_1_sva(1)) XOR (input_sva(59)) XOR (s_output_1_19_16_50_sva(3)));
  s_output_1_3_0_40_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_19_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_23_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_23_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_23_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_23_rg_addr <= STD_LOGIC_VECTOR'( "111")
      & ((input_sva(25)) XOR (s_output_1_19_16_35_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(42)))
      & ((input_sva(7)) XOR (s_output_1_19_16_5_sva(0)) XOR (key_io_read_key_rsc_cse_63_1_sva(56)))
      & ((input_sva(33)) XOR (s_output_1_3_0_39_sva(2)) XOR (key_io_read_key_rsc_cse_63_1_sva(10)))
      & ((input_sva(41)) XOR (s_output_1_19_16_50_sva(1)) XOR (key_io_read_key_rsc_cse_63_1_sva(43)))
      & ((input_sva(49)) XOR (s_output_1_19_16_20_sva(0)) XOR (key_io_read_key_rsc_cse_63_1_sva(25)))
      & ((input_sva(57)) XOR (s_output_1_3_0_54_sva(3)) XOR (key_io_read_key_rsc_cse_63_1_sva(32)));
  s_output_1_3_0_10_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_23_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_30_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_30_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_30_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_30_rg_addr <= STD_LOGIC_VECTOR'( "011")
      & (R_20_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(44))) & (R_15_3_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(62))) & (R_19_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(37)))
      & (R_18_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(38))) & (R_17_3_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(11))) & (R_16_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(20)));
  s_output_1_19_16_7_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_30_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_29_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_29_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_29_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_29_rg_addr <= STD_LOGIC_VECTOR'( "110")
      & (R_8_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(42))) & (R_3_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(16)))
      & (R_7_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(51))) & (R_6_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(2)))
      & (R_5_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(40))) & (R_4_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(25)));
  s_output_1_3_0_56_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_29_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_26_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_26_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_26_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_26_rg_addr <= STD_LOGIC_VECTOR'( "001")
      & (R_28_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(5))) & (R_23_3_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(61))) & (R_27_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(46)))
      & (R_26_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(36))) & (R_25_3_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(29))) & (R_24_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(19)));
  s_output_1_19_16_37_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_26_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_24_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_24_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_24_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_24_rg_addr <= STD_LOGIC_VECTOR'( "000")
      & (R_0_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(28))) & (R_27_3_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(21))) & (R_31_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(52)))
      & (R_30_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(4))) & (R_29_3_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(14))) & (R_28_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(54)));
  s_output_1_19_16_22_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_24_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_25_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_25_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_25_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_25_rg_addr <= STD_LOGIC_VECTOR'( "100")
      & (R_16_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(18))) & (R_11_3_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(32))) & (R_15_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(8)))
      & (R_14_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(1))) & (R_13_3_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(49))) & (R_12_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(35)));
  s_output_1_3_0_26_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_25_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_28_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_28_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_28_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_28_rg_addr <= STD_LOGIC_VECTOR'( "010")
      & (R_24_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(6))) & (R_19_3_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(45))) & (R_23_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(3)))
      & (R_22_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(12))) & (R_21_3_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(13))) & (R_20_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(30)));
  s_output_1_19_16_52_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_28_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_27_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_27_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_27_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_27_rg_addr <= STD_LOGIC_VECTOR'( "101")
      & (R_12_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(56))) & (R_7_3_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(43))) & (R_11_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(10)))
      & (R_10_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(0))) & (R_9_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(50)))
      & (R_8_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(17)));
  s_output_1_3_0_41_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_27_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_31_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_31_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_31_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_31_rg_addr <= STD_LOGIC_VECTOR'( "111")
      & (R_4_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(58))) & (R_31_3_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(9))) & (R_3_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(26)))
      & (R_2_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(59))) & (R_1_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(41)))
      & (R_0_3_sva XOR (key_io_read_key_rsc_cse_63_1_sva(48)));
  s_output_1_3_0_11_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_31_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_38_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_38_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_38_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_38_rg_addr <= STD_LOGIC_VECTOR'( "011")
      & (R_20_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(60))) & (R_15_4_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(13))) & (R_19_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(53)))
      & (R_18_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(54))) & (R_17_4_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(27))) & (R_16_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(36)));
  s_output_1_19_16_8_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_38_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_37_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_37_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_37_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_37_rg_addr <= STD_LOGIC_VECTOR'( "110")
      & (R_8_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(58))) & (R_3_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(32)))
      & (R_7_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(0))) & (R_6_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(18)))
      & (R_5_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(56))) & (R_4_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(41)));
  s_output_1_3_0_57_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_37_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_34_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_34_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_34_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_34_rg_addr <= STD_LOGIC_VECTOR'( "001")
      & (R_28_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(21))) & (R_23_4_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(12))) & (R_27_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(62)))
      & (R_26_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(52))) & (R_25_4_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(45))) & (R_24_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(6)));
  s_output_1_19_16_38_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_34_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_32_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_32_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_32_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_32_rg_addr <= STD_LOGIC_VECTOR'( "000")
      & (R_0_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(44))) & (R_27_4_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(37))) & (R_31_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(3)))
      & (R_30_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(20))) & (R_29_4_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(30))) & (R_28_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(5)));
  s_output_1_19_16_23_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_32_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_33_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_33_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_33_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_33_rg_addr <= STD_LOGIC_VECTOR'( "100")
      & (R_16_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(34))) & (R_11_4_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(48))) & (R_15_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(24)))
      & (R_14_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(17))) & (R_13_4_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(2))) & (R_12_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(51)));
  s_output_1_3_0_27_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_33_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_36_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_36_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_36_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_36_rg_addr <= STD_LOGIC_VECTOR'( "010")
      & (R_24_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(22))) & (R_19_4_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(61))) & (R_23_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(19)))
      & (R_22_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(28))) & (R_21_4_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(29))) & (R_20_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(46)));
  s_output_1_19_16_53_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_36_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_35_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_35_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_35_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_35_rg_addr <= STD_LOGIC_VECTOR'( "101")
      & (R_12_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(9))) & (R_7_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(59)))
      & (R_11_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(26))) & (R_10_4_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(16))) & (R_9_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(35)))
      & (R_8_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(33)));
  s_output_1_3_0_42_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_35_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_39_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_39_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_39_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_39_rg_addr <= STD_LOGIC_VECTOR'( "111")
      & (R_4_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(43))) & (R_31_4_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(25))) & (R_3_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(42)))
      & (R_2_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(8))) & (R_1_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(57)))
      & (R_0_4_sva XOR (key_io_read_key_rsc_cse_63_1_sva(1)));
  s_output_1_3_0_12_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_39_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_46_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_46_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_46_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_46_rg_addr <= STD_LOGIC_VECTOR'( "011")
      & (R_20_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(11))) & (R_15_5_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(29))) & (R_19_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(4)))
      & (R_18_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(5))) & (R_17_5_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(14))) & (R_16_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(52)));
  s_output_1_19_16_9_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_46_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_45_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_45_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_45_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_45_rg_addr <= STD_LOGIC_VECTOR'( "110")
      & (R_8_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(43))) & (R_3_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(48)))
      & (R_7_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(16))) & (R_6_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(34)))
      & (R_5_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(9))) & (R_4_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(57)));
  s_output_1_3_0_58_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_45_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_42_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_42_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_42_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_42_rg_addr <= STD_LOGIC_VECTOR'( "001")
      & (R_28_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(37))) & (R_23_5_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(28))) & (R_27_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(13)))
      & (R_26_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(3))) & (R_25_5_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(61))) & (R_24_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(22)));
  s_output_1_19_16_39_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_42_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_40_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_40_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_40_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_40_rg_addr <= STD_LOGIC_VECTOR'( "000")
      & (R_0_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(60))) & (R_27_5_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(53))) & (R_31_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(19)))
      & (R_30_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(36))) & (R_29_5_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(46))) & (R_28_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(21)));
  s_output_1_19_16_24_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_40_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_41_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_41_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_41_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_41_rg_addr <= STD_LOGIC_VECTOR'( "100")
      & (R_16_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(50))) & (R_11_5_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(1))) & (R_15_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(40)))
      & (R_14_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(33))) & (R_13_5_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(18))) & (R_12_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(0)));
  s_output_1_3_0_28_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_41_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_44_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_44_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_44_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_44_rg_addr <= STD_LOGIC_VECTOR'( "010")
      & (R_24_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(38))) & (R_19_5_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(12))) & (R_23_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(6)))
      & (R_22_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(44))) & (R_21_5_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(45))) & (R_20_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(62)));
  s_output_1_19_16_54_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_44_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_43_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_43_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_43_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_43_rg_addr <= STD_LOGIC_VECTOR'( "101")
      & (R_12_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(25))) & (R_7_5_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(8))) & (R_11_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(42)))
      & (R_10_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(32))) & (R_9_5_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(51))) & (R_8_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(49)));
  s_output_1_3_0_43_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_43_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_47_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_47_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_47_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_47_rg_addr <= STD_LOGIC_VECTOR'( "111")
      & (R_4_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(59))) & (R_31_5_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(41))) & (R_3_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(58)))
      & (R_2_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(24))) & (R_1_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(10)))
      & (R_0_5_sva XOR (key_io_read_key_rsc_cse_63_1_sva(17)));
  s_output_1_3_0_13_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_47_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_54_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_54_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_54_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_54_rg_addr <= STD_LOGIC_VECTOR'( "011")
      & (R_20_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(27))) & (R_15_6_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(45))) & (R_19_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(20)))
      & (R_18_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(21))) & (R_17_6_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(30))) & (R_16_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(3)));
  s_output_1_19_16_10_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_54_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_53_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_53_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_53_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_53_rg_addr <= STD_LOGIC_VECTOR'( "110")
      & (R_8_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(59))) & (R_3_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(1)))
      & (R_7_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(32))) & (R_6_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(50)))
      & (R_5_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(25))) & (R_4_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(10)));
  s_output_1_3_0_59_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_53_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_50_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_50_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_50_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_50_rg_addr <= STD_LOGIC_VECTOR'( "001")
      & (R_28_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(53))) & (R_23_6_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(44))) & (R_27_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(29)))
      & (R_26_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(19))) & (R_25_6_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(12))) & (R_24_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(38)));
  s_output_1_19_16_40_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_50_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_48_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_48_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_48_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_48_rg_addr <= STD_LOGIC_VECTOR'( "000")
      & (R_0_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(11))) & (R_27_6_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(4))) & (R_31_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(6)))
      & (R_30_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(52))) & (R_29_6_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(62))) & (R_28_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(37)));
  s_output_1_19_16_25_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_48_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_49_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_49_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_49_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_49_rg_addr <= STD_LOGIC_VECTOR'( "100")
      & (R_16_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(35))) & (R_11_6_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(17))) & (R_15_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(56)))
      & (R_14_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(49))) & (R_13_6_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(34))) & (R_12_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(16)));
  s_output_1_3_0_29_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_49_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_52_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_52_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_52_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_52_rg_addr <= STD_LOGIC_VECTOR'( "010")
      & (R_24_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(54))) & (R_19_6_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(28))) & (R_23_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(22)))
      & (R_22_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(60))) & (R_21_6_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(61))) & (R_20_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(13)));
  s_output_1_19_16_55_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_52_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_51_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_51_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_51_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_51_rg_addr <= STD_LOGIC_VECTOR'( "101")
      & (R_12_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(41))) & (R_7_6_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(24))) & (R_11_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(58)))
      & (R_10_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(48))) & (R_9_6_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(0))) & (R_8_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(2)));
  s_output_1_3_0_44_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_51_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_55_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_55_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_55_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_55_rg_addr <= STD_LOGIC_VECTOR'( "111")
      & (R_4_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(8))) & (R_31_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(57)))
      & (R_3_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(43))) & (R_2_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(40)))
      & (R_1_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(26))) & (R_0_6_sva XOR (key_io_read_key_rsc_cse_63_1_sva(33)));
  s_output_1_3_0_14_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_55_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_62_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_62_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_62_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_62_rg_addr <= STD_LOGIC_VECTOR'( "011")
      & (R_20_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(14))) & (R_15_7_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(61))) & (R_19_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(36)))
      & (R_18_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(37))) & (R_17_7_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(46))) & (R_16_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(19)));
  s_output_1_19_16_11_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_62_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_61_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_61_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_61_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_61_rg_addr <= STD_LOGIC_VECTOR'( "110")
      & (R_8_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(8))) & (R_3_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(17)))
      & (R_7_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(48))) & (R_6_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(35)))
      & (R_5_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(41))) & (R_4_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(26)));
  s_output_1_3_0_60_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_61_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_58_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_58_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_58_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_58_rg_addr <= STD_LOGIC_VECTOR'( "001")
      & (R_28_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(4))) & (R_23_7_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(60))) & (R_27_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(45)))
      & (R_26_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(6))) & (R_25_7_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(28))) & (R_24_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(54)));
  s_output_1_19_16_41_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_58_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_56_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_56_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_56_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_56_rg_addr <= STD_LOGIC_VECTOR'( "000")
      & (R_0_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(27))) & (R_27_7_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(20))) & (R_31_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(22)))
      & (R_30_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(3))) & (R_29_7_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(13))) & (R_28_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(53)));
  s_output_1_19_16_26_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_56_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_57_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_57_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_57_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_57_rg_addr <= STD_LOGIC_VECTOR'( "100")
      & (R_16_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(51))) & (R_11_7_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(33))) & (R_15_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(9)))
      & (R_14_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(2))) & (R_13_7_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(50))) & (R_12_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(32)));
  s_output_1_3_0_30_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_57_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_60_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_60_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_60_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_60_rg_addr <= STD_LOGIC_VECTOR'( "010")
      & (R_24_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(5))) & (R_19_7_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(44))) & (R_23_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(38)))
      & (R_22_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(11))) & (R_21_7_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(12))) & (R_20_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(29)));
  s_output_1_19_16_56_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_60_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_59_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_59_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_59_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_59_rg_addr <= STD_LOGIC_VECTOR'( "101")
      & (R_12_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(57))) & (R_7_7_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(40))) & (R_11_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(43)))
      & (R_10_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(1))) & (R_9_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(16)))
      & (R_8_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(18)));
  s_output_1_3_0_45_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_59_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_63_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_63_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_63_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_63_rg_addr <= STD_LOGIC_VECTOR'( "111")
      & (R_4_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(24))) & (R_31_7_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(10))) & (R_3_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(59)))
      & (R_2_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(56))) & (R_1_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(42)))
      & (R_0_7_sva XOR (key_io_read_key_rsc_cse_63_1_sva(49)));
  s_output_1_3_0_15_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_63_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_70_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_70_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_70_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_70_rg_addr <= STD_LOGIC_VECTOR'( "011")
      & (R_20_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(22))) & (R_15_8_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(4))) & (R_19_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(44)))
      & (R_18_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(45))) & (R_17_8_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(54))) & (R_16_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(27)));
  s_output_1_19_16_12_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_70_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_69_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_69_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_69_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_69_rg_addr <= STD_LOGIC_VECTOR'( "110")
      & (R_8_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(16))) & (R_3_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(25)))
      & (R_7_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(56))) & (R_6_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(43)))
      & (R_5_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(49))) & (R_4_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(34)));
  s_output_1_3_0_61_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_69_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_66_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_66_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_66_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_66_rg_addr <= STD_LOGIC_VECTOR'( "001")
      & (R_28_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(12))) & (R_23_8_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(3))) & (R_27_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(53)))
      & (R_26_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(14))) & (R_25_8_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(36))) & (R_24_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(62)));
  s_output_1_19_16_42_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_66_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_64_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_64_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_64_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_64_rg_addr <= STD_LOGIC_VECTOR'( "000")
      & (R_0_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(6))) & (R_27_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(28)))
      & (R_31_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(30))) & (R_30_8_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(11))) & (R_29_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(21)))
      & (R_28_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(61)));
  s_output_1_19_16_27_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_64_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_65_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_65_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_65_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_65_rg_addr <= STD_LOGIC_VECTOR'( "100")
      & (R_16_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(59))) & (R_11_8_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(41))) & (R_15_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(17)))
      & (R_14_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(10))) & (R_13_8_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(58))) & (R_12_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(40)));
  s_output_1_3_0_31_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_65_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_68_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_68_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_68_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_68_rg_addr <= STD_LOGIC_VECTOR'( "010")
      & (R_24_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(13))) & (R_19_8_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(52))) & (R_23_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(46)))
      & (R_22_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(19))) & (R_21_8_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(20))) & (R_20_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(37)));
  s_output_1_19_16_57_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_68_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_67_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_67_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_67_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_67_rg_addr <= STD_LOGIC_VECTOR'( "101")
      & (R_12_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(2))) & (R_7_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(48)))
      & (R_11_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(51))) & (R_10_8_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(9))) & (R_9_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(24)))
      & (R_8_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(26)));
  s_output_1_3_0_46_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_67_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_71_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_71_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_71_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_71_rg_addr <= STD_LOGIC_VECTOR'( "111")
      & (R_4_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(32))) & (R_31_8_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(18))) & (R_3_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(0)))
      & (R_2_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(1))) & (R_1_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(50)))
      & (R_0_8_sva XOR (key_io_read_key_rsc_cse_63_1_sva(57)));
  s_output_1_3_0_16_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_71_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_78_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_78_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_78_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_78_rg_addr <= STD_LOGIC_VECTOR'( "011")
      & (R_20_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(38))) & (R_15_9_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(20))) & (R_19_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(60)))
      & (R_18_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(61))) & (R_17_9_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(5))) & (R_16_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(14)));
  s_output_1_19_16_13_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_78_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_77_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_77_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_77_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_77_rg_addr <= STD_LOGIC_VECTOR'( "110")
      & (R_8_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(32))) & (R_3_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(41)))
      & (R_7_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(9))) & (R_6_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(59)))
      & (R_5_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(2))) & (R_4_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(50)));
  s_output_1_3_0_62_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_77_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_74_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_74_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_74_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_74_rg_addr <= STD_LOGIC_VECTOR'( "001")
      & (R_28_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(28))) & (R_23_9_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(19))) & (R_27_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(4)))
      & (R_26_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(30))) & (R_25_9_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(52))) & (R_24_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(13)));
  s_output_1_19_16_43_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_74_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_72_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_72_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_72_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_72_rg_addr <= STD_LOGIC_VECTOR'( "000")
      & (R_0_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(22))) & (R_27_9_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(44))) & (R_31_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(46)))
      & (R_30_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(27))) & (R_29_9_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(37))) & (R_28_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(12)));
  s_output_1_19_16_28_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_72_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_73_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_73_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_73_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_73_rg_addr <= STD_LOGIC_VECTOR'( "100")
      & (R_16_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(8))) & (R_11_9_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(57))) & (R_15_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(33)))
      & (R_14_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(26))) & (R_13_9_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(43))) & (R_12_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(56)));
  s_output_1_3_0_32_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_73_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_76_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_76_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_76_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_76_rg_addr <= STD_LOGIC_VECTOR'( "010")
      & (R_24_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(29))) & (R_19_9_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(3))) & (R_23_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(62)))
      & (R_22_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(6))) & (R_21_9_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(36))) & (R_20_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(53)));
  s_output_1_19_16_58_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_76_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_75_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_75_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_75_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_75_rg_addr <= STD_LOGIC_VECTOR'( "101")
      & (R_12_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(18))) & (R_7_9_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(1))) & (R_11_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(0)))
      & (R_10_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(25))) & (R_9_9_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(40))) & (R_8_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(42)));
  s_output_1_3_0_47_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_75_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_79_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_79_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_79_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_79_rg_addr <= STD_LOGIC_VECTOR'( "111")
      & (R_4_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(48))) & (R_31_9_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(34))) & (R_3_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(16)))
      & (R_2_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(17))) & (R_1_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(35)))
      & (R_0_9_sva XOR (key_io_read_key_rsc_cse_63_1_sva(10)));
  s_output_1_3_0_17_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_79_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_86_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_86_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_86_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_86_rg_addr <= STD_LOGIC_VECTOR'( "011")
      & (R_20_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(54))) & (R_15_10_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(36))) & (R_19_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(11)))
      & (R_18_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(12))) & (R_17_10_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(21))) & (R_16_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(30)));
  s_output_1_19_16_14_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_86_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_85_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_85_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_85_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_85_rg_addr <= STD_LOGIC_VECTOR'( "110")
      & (R_8_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(48))) & (R_3_10_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(57))) & (R_7_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(25)))
      & (R_6_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(8))) & (R_5_10_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(18))) & (R_4_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(35)));
  s_output_1_3_0_63_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_85_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_82_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_82_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_82_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_82_rg_addr <= STD_LOGIC_VECTOR'( "001")
      & (R_28_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(44))) & (R_23_10_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(6))) & (R_27_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(20)))
      & (R_26_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(46))) & (R_25_10_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(3))) & (R_24_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(29)));
  s_output_1_19_16_44_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_82_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_80_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_80_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_80_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_80_rg_addr <= STD_LOGIC_VECTOR'( "000")
      & (R_0_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(38))) & (R_27_10_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(60))) & (R_31_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(62)))
      & (R_30_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(14))) & (R_29_10_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(53))) & (R_28_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(28)));
  s_output_1_19_16_29_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_80_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_81_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_81_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_81_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_81_rg_addr <= STD_LOGIC_VECTOR'( "100")
      & (R_16_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(24))) & (R_11_10_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(10))) & (R_15_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(49)))
      & (R_14_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(42))) & (R_13_10_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(59))) & (R_12_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(9)));
  s_output_1_3_0_33_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_81_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_84_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_84_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_84_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_84_rg_addr <= STD_LOGIC_VECTOR'( "010")
      & (R_24_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(45))) & (R_19_10_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(19))) & (R_23_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(13)))
      & (R_22_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(22))) & (R_21_10_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(52))) & (R_20_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(4)));
  s_output_1_19_16_59_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_84_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_83_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_83_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_83_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_83_rg_addr <= STD_LOGIC_VECTOR'( "101")
      & (R_12_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(34))) & (R_7_10_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(17))) & (R_11_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(16)))
      & (R_10_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(41))) & (R_9_10_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(56))) & (R_8_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(58)));
  s_output_1_3_0_48_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_83_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_87_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_87_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_87_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_87_rg_addr <= STD_LOGIC_VECTOR'( "111")
      & (R_4_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(1))) & (R_31_10_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(50))) & (R_3_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(32)))
      & (R_2_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(33))) & (R_1_10_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(51))) & (R_0_10_sva XOR (key_io_read_key_rsc_cse_63_1_sva(26)));
  s_output_1_3_0_18_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_87_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_94_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_94_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_94_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_94_rg_addr <= STD_LOGIC_VECTOR'( "011")
      & (R_20_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(5))) & (R_15_11_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(52))) & (R_19_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(27)))
      & (R_18_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(28))) & (R_17_11_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(37))) & (R_16_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(46)));
  s_output_1_19_16_15_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_94_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_93_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_93_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_93_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_93_rg_addr <= STD_LOGIC_VECTOR'( "110")
      & (R_8_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(1))) & (R_3_11_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(10))) & (R_7_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(41)))
      & (R_6_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(24))) & (R_5_11_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(34))) & (R_4_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(51)));
  s_output_1_3_0_64_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_93_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_90_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_90_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_90_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_90_rg_addr <= STD_LOGIC_VECTOR'( "001")
      & (R_28_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(60))) & (R_23_11_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(22))) & (R_27_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(36)))
      & (R_26_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(62))) & (R_25_11_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(19))) & (R_24_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(45)));
  s_output_1_19_16_45_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_90_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_88_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_88_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_88_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_88_rg_addr <= STD_LOGIC_VECTOR'( "000")
      & (R_0_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(54))) & (R_27_11_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(11))) & (R_31_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(13)))
      & (R_30_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(30))) & (R_29_11_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(4))) & (R_28_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(44)));
  s_output_1_19_16_30_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_88_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_89_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_89_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_89_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_89_rg_addr <= STD_LOGIC_VECTOR'( "100")
      & (R_16_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(40))) & (R_11_11_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(26))) & (R_15_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(2)))
      & (R_14_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(58))) & (R_13_11_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(8))) & (R_12_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(25)));
  s_output_1_3_0_34_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_89_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_92_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_92_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_92_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_92_rg_addr <= STD_LOGIC_VECTOR'( "010")
      & (R_24_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(61))) & (R_19_11_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(6))) & (R_23_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(29)))
      & (R_22_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(38))) & (R_21_11_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(3))) & (R_20_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(20)));
  s_output_1_19_16_60_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_92_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_91_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_91_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_91_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_91_rg_addr <= STD_LOGIC_VECTOR'( "101")
      & (R_12_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(50))) & (R_7_11_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(33))) & (R_11_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(32)))
      & (R_10_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(57))) & (R_9_11_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(9))) & (R_8_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(43)));
  s_output_1_3_0_49_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_91_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_95_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_95_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_95_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_95_rg_addr <= STD_LOGIC_VECTOR'( "111")
      & (R_4_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(17))) & (R_31_11_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(35))) & (R_3_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(48)))
      & (R_2_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(49))) & (R_1_11_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(0))) & (R_0_11_sva XOR (key_io_read_key_rsc_cse_63_1_sva(42)));
  s_output_1_3_0_19_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_95_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_102_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_102_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_102_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_102_rg_addr <= STD_LOGIC_VECTOR'( "011")
      & (R_20_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(21))) & (R_15_12_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(3))) & (R_19_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(14)))
      & (R_18_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(44))) & (R_17_12_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(53))) & (R_16_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(62)));
  s_output_1_19_16_16_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_102_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_101_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_101_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_101_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_101_rg_addr <= STD_LOGIC_VECTOR'( "110")
      & (R_8_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(17))) & (R_3_12_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(26))) & (R_7_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(57)))
      & (R_6_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(40))) & (R_5_12_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(50))) & (R_4_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(0)));
  s_output_1_3_0_65_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_101_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_98_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_98_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_98_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_98_rg_addr <= STD_LOGIC_VECTOR'( "001")
      & (R_28_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(11))) & (R_23_12_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(38))) & (R_27_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(52)))
      & (R_26_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(13))) & (R_25_12_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(6))) & (R_24_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(61)));
  s_output_1_19_16_46_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_98_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_96_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_96_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_96_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_96_rg_addr <= STD_LOGIC_VECTOR'( "000")
      & (R_0_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(5))) & (R_27_12_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(27))) & (R_31_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(29)))
      & (R_30_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(46))) & (R_29_12_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(20))) & (R_28_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(60)));
  s_output_1_19_16_31_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_96_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_97_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_97_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_97_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_97_rg_addr <= STD_LOGIC_VECTOR'( "100")
      & (R_16_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(56))) & (R_11_12_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(42))) & (R_15_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(18)))
      & (R_14_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(43))) & (R_13_12_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(24))) & (R_12_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(41)));
  s_output_1_3_0_35_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_97_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_100_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_100_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_100_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_100_rg_addr <= STD_LOGIC_VECTOR'( "010")
      & (R_24_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(12))) & (R_19_12_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(22))) & (R_23_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(45)))
      & (R_22_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(54))) & (R_21_12_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(19))) & (R_20_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(36)));
  s_output_1_19_16_61_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_100_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_99_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_99_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_99_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_99_rg_addr <= STD_LOGIC_VECTOR'( "101")
      & (R_12_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(35))) & (R_7_12_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(49))) & (R_11_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(48)))
      & (R_10_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(10))) & (R_9_12_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(25))) & (R_8_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(59)));
  s_output_1_3_0_50_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_99_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_103_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_103_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_103_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_103_rg_addr <= STD_LOGIC_VECTOR'( "111")
      & (R_4_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(33))) & (R_31_12_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(51))) & (R_3_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(1)))
      & (R_2_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(2))) & (R_1_12_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(16))) & (R_0_12_sva XOR (key_io_read_key_rsc_cse_63_1_sva(58)));
  s_output_1_3_0_20_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_103_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_110_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_110_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_110_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_110_rg_addr <= STD_LOGIC_VECTOR'( "011")
      & (R_20_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(37))) & (R_15_13_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(19))) & (R_19_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(30)))
      & (R_18_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(60))) & (R_17_13_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(4))) & (R_16_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(13)));
  s_output_1_19_16_17_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_110_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_109_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_109_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_109_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_109_rg_addr <= STD_LOGIC_VECTOR'( "110")
      & (R_8_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(33))) & (R_3_13_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(42))) & (R_7_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(10)))
      & (R_6_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(56))) & (R_5_13_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(35))) & (R_4_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(16)));
  s_output_1_3_0_66_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_109_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_106_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_106_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_106_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_106_rg_addr <= STD_LOGIC_VECTOR'( "001")
      & (R_28_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(27))) & (R_23_13_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(54))) & (R_27_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(3)))
      & (R_26_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(29))) & (R_25_13_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(22))) & (R_24_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(12)));
  s_output_1_19_16_47_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_106_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_104_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_104_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_104_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_104_rg_addr <= STD_LOGIC_VECTOR'( "000")
      & (R_0_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(21))) & (R_27_13_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(14))) & (R_31_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(45)))
      & (R_30_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(62))) & (R_29_13_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(36))) & (R_28_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(11)));
  s_output_1_19_16_32_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_104_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_105_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_105_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_105_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_105_rg_addr <= STD_LOGIC_VECTOR'( "100")
      & (R_16_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(9))) & (R_11_13_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(58))) & (R_15_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(34)))
      & (R_14_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(59))) & (R_13_13_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(40))) & (R_12_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(57)));
  s_output_1_3_0_36_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_105_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_108_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_108_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_108_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_108_rg_addr <= STD_LOGIC_VECTOR'( "010")
      & (R_24_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(28))) & (R_19_13_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(38))) & (R_23_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(61)))
      & (R_22_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(5))) & (R_21_13_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(6))) & (R_20_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(52)));
  s_output_1_19_16_62_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_108_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_107_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_107_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_107_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_107_rg_addr <= STD_LOGIC_VECTOR'( "101")
      & (R_12_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(51))) & (R_7_13_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(2))) & (R_11_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(1)))
      & (R_10_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(26))) & (R_9_13_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(41))) & (R_8_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(8)));
  s_output_1_3_0_51_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_107_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_111_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_111_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_111_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_111_rg_addr <= STD_LOGIC_VECTOR'( "111")
      & (R_4_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(49))) & (R_31_13_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(0))) & (R_3_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(17)))
      & (R_2_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(18))) & (R_1_13_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(32))) & (R_0_13_sva XOR (key_io_read_key_rsc_cse_63_1_sva(43)));
  s_output_1_3_0_21_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_111_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_118_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_118_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_118_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_118_rg_addr <= STD_LOGIC_VECTOR'( "011")
      & (R_20_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(53))) & (R_15_14_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(6))) & (R_19_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(46)))
      & (R_18_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(11))) & (R_17_14_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(20))) & (R_16_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(29)));
  s_output_1_19_16_18_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_118_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_117_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_117_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_117_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_117_rg_addr <= STD_LOGIC_VECTOR'( "110")
      & (R_8_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(49))) & (R_3_14_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(58))) & (R_7_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(26)))
      & (R_6_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(9))) & (R_5_14_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(51))) & (R_4_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(32)));
  s_output_1_3_0_67_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_117_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_114_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_114_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_114_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_114_rg_addr <= STD_LOGIC_VECTOR'( "001")
      & (R_28_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(14))) & (R_23_14_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(5))) & (R_27_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(19)))
      & (R_26_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(45))) & (R_25_14_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(38))) & (R_24_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(28)));
  s_output_1_19_16_48_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_114_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_112_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_112_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_112_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_112_rg_addr <= STD_LOGIC_VECTOR'( "000")
      & (R_0_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(37))) & (R_27_14_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(30))) & (R_31_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(61)))
      & (R_30_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(13))) & (R_29_14_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(52))) & (R_28_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(27)));
  s_output_1_19_16_33_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_112_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_113_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_113_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_113_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_113_rg_addr <= STD_LOGIC_VECTOR'( "100")
      & (R_16_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(25))) & (R_11_14_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(43))) & (R_15_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(50)))
      & (R_14_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(8))) & (R_13_14_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(56))) & (R_12_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(10)));
  s_output_1_3_0_37_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_113_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_116_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_116_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_116_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_116_rg_addr <= STD_LOGIC_VECTOR'( "010")
      & (R_24_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(44))) & (R_19_14_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(54))) & (R_23_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(12)))
      & (R_22_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(21))) & (R_21_14_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(22))) & (R_20_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(3)));
  s_output_1_19_16_63_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_116_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_115_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_115_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_115_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_115_rg_addr <= STD_LOGIC_VECTOR'( "101")
      & (R_12_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(0))) & (R_7_14_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(18))) & (R_11_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(17)))
      & (R_10_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(42))) & (R_9_14_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(57))) & (R_8_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(24)));
  s_output_1_3_0_52_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_115_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_119_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_119_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_119_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_119_rg_addr <= STD_LOGIC_VECTOR'( "111")
      & (R_4_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(2))) & (R_31_14_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(16))) & (R_3_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(33)))
      & (R_2_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(34))) & (R_1_14_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(48))) & (R_0_14_sva XOR (key_io_read_key_rsc_cse_63_1_sva(59)));
  s_output_1_3_0_22_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_119_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_121_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_121_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_121_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_121_rg_addr <= STD_LOGIC_VECTOR'( "100")
      & (R_16_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(33))) & (R_11_15_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(51))) & (R_15_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(58)))
      & (R_14_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(16))) & (R_13_15_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(1))) & (R_12_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(18)));
  s_output_1_3_0_5_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_121_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_120_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_120_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_120_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_120_rg_addr <= STD_LOGIC_VECTOR'( "000")
      & (R_0_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(45))) & (R_27_15_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(38))) & (R_31_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(4)))
      & (R_30_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(21))) & (R_29_15_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(60))) & (R_28_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(6)));
  s_output_1_19_16_1_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_120_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_124_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_124_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_124_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_124_rg_addr <= STD_LOGIC_VECTOR'( "010")
      & (R_24_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(52))) & (R_19_15_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(62))) & (R_23_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(20)))
      & (R_22_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(29))) & (R_21_15_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(30))) & (R_20_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(11)));
  s_output_1_19_16_3_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_124_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_126_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_126_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_126_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_126_rg_addr <= STD_LOGIC_VECTOR'( "011")
      & (R_20_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(61))) & (R_15_15_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(14))) & (R_19_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(54)))
      & (R_18_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(19))) & (R_17_15_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(28))) & (R_16_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(37)));
  s_output_1_19_16_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_126_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_125_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_125_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_125_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_125_rg_addr <= STD_LOGIC_VECTOR'( "110")
      & (R_8_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(57))) & (R_3_15_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(35))) & (R_7_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(34)))
      & (R_6_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(17))) & (R_5_15_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(59))) & (R_4_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(40)));
  s_output_1_3_0_7_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_125_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_122_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_122_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_122_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_122_rg_addr <= STD_LOGIC_VECTOR'( "001")
      & (R_28_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(22))) & (R_23_15_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(13))) & (R_27_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(27)))
      & (R_26_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(53))) & (R_25_15_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(46))) & (R_24_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(36)));
  s_output_1_19_16_2_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_122_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_127_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_127_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_127_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_127_rg_addr <= STD_LOGIC_VECTOR'( "111")
      & (R_4_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(10))) & (R_31_15_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(24))) & (R_3_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(41)))
      & (R_2_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(42))) & (R_1_15_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(56))) & (R_0_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(0)));
  s_output_1_3_0_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_127_rg_data_out;

  operator_8_false_1_read_rom_S_rom_map_1_123_rg : work.des_checkmgc_rom_12_512_4_1_pkg.des_checkmgc_rom_12_512_4_1
    PORT MAP(
      addr => operator_8_false_1_read_rom_S_rom_map_1_123_rg_addr,
      data_out => operator_8_false_1_read_rom_S_rom_map_1_123_rg_data_out
    );
  operator_8_false_1_read_rom_S_rom_map_1_123_rg_addr <= STD_LOGIC_VECTOR'( "101")
      & (R_12_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(8))) & (R_7_15_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(26))) & (R_11_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(25)))
      & (R_10_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(50))) & (R_9_15_sva XOR
      (key_io_read_key_rsc_cse_63_1_sva(2))) & (R_8_15_sva XOR (key_io_read_key_rsc_cse_63_1_sva(32)));
  s_output_1_3_0_6_sva_1 <= operator_8_false_1_read_rom_S_rom_map_1_123_rg_data_out;

  des_check_core_core_fsm_inst : des_check_core_core_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      fsm_output => des_check_core_core_fsm_inst_fsm_output
    );
  fsm_output <= des_check_core_core_fsm_inst_fsm_output;

  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(0)) = '1' ) THEN
        key_io_read_key_rsc_cse_63_1_sva <= key_rsci_idat(63 DOWNTO 1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_31 <= R_28_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_32 <= R_3_14_sva XOR (s_output_1_3_0_6_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_30 <= R_28_14_sva XOR (s_output_1_3_0_6_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_33 <= R_3_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_29 <= R_20_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_34 <= R_11_14_sva XOR (s_output_1_3_0_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_28 <= R_20_14_sva XOR (s_output_1_3_0_7_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_35 <= R_11_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_27 <= R_12_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_36 <= R_19_14_sva XOR (s_output_1_19_16_2_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_26 <= R_12_14_sva XOR (s_output_1_19_16_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_37 <= R_19_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_25 <= R_4_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_38 <= R_27_14_sva XOR (s_output_1_3_0_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_24 <= R_4_14_sva XOR (s_output_1_19_16_2_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_39 <= R_27_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_23 <= R_29_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_40 <= R_2_14_sva XOR (s_output_1_19_16_3_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_22 <= R_29_14_sva XOR (s_output_1_3_0_5_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_41 <= R_2_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_21 <= R_21_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_42 <= R_10_14_sva XOR (s_output_1_3_0_7_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_20 <= R_21_14_sva XOR (s_output_1_3_0_6_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_43 <= R_10_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_19 <= R_13_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_44 <= R_18_14_sva XOR (s_output_1_3_0_5_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_18 <= R_13_14_sva XOR (s_output_1_3_0_6_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_45 <= R_18_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_17 <= R_5_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_46 <= R_26_14_sva XOR (s_output_1_19_16_3_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_16 <= R_5_14_sva XOR (s_output_1_3_0_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_47 <= R_26_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_15 <= R_30_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_48 <= R_1_14_sva XOR (s_output_1_19_16_1_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_14 <= R_30_14_sva XOR (s_output_1_19_16_2_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_49 <= R_1_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_13 <= R_22_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_50 <= R_9_14_sva XOR (s_output_1_19_16_1_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_12 <= R_22_14_sva XOR (s_output_1_19_16_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_51 <= R_9_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_11 <= R_14_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_52 <= R_17_14_sva XOR (s_output_1_3_0_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_10 <= R_14_14_sva XOR (s_output_1_19_16_2_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_53 <= R_17_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_9 <= R_6_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_54 <= R_25_14_sva XOR (s_output_1_3_0_7_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_8 <= R_6_14_sva XOR (s_output_1_19_16_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_55 <= R_25_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_7 <= R_31_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_56 <= R_0_14_sva XOR (s_output_1_3_0_7_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_6 <= R_31_14_sva XOR (s_output_1_19_16_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_57 <= R_0_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_5 <= R_23_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_58 <= R_8_14_sva XOR (s_output_1_19_16_3_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_4 <= R_23_14_sva XOR (s_output_1_19_16_1_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_59 <= R_8_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_3 <= R_15_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_60 <= R_16_14_sva XOR (s_output_1_19_16_3_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_2 <= R_15_14_sva XOR (s_output_1_19_16_1_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_61 <= R_16_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_1 <= R_7_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_62 <= R_24_14_sva XOR (s_output_1_3_0_5_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_0 <= R_7_14_sva XOR (s_output_1_3_0_5_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(15)) = '1' ) THEN
        return_rsci_idat_63 <= R_24_15_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(0)) = '1' ) THEN
        input_sva <= input_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_input_rsc_triosy_obj_ld_cse <= '0';
        return_rsc_triosy_obj_ld <= '0';
      ELSE
        reg_input_rsc_triosy_obj_ld_cse <= fsm_output(0);
        return_rsc_triosy_obj_ld <= fsm_output(15);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      s_output_1_19_16_4_sva <= operator_8_false_1_read_rom_S_rom_map_1_6_itm;
      s_output_1_3_0_53_sva <= operator_8_false_1_read_rom_S_rom_map_1_5_itm;
      s_output_1_19_16_34_sva <= operator_8_false_1_read_rom_S_rom_map_1_2_itm;
      s_output_1_19_16_19_sva <= operator_8_false_1_read_rom_S_rom_map_1_itm;
      s_output_1_3_0_23_sva <= operator_8_false_1_read_rom_S_rom_map_1_1_itm;
      s_output_1_19_16_49_sva <= operator_8_false_1_read_rom_S_rom_map_1_4_itm;
      s_output_1_3_0_38_sva <= operator_8_false_1_read_rom_S_rom_map_1_3_itm;
      s_output_1_3_0_8_sva <= operator_8_false_1_read_rom_S_rom_map_1_7_itm;
      R_31_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_32_nl, loop_DES_rounds_2_xor_32_nl,
          fsm_output(2));
      R_0_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_31_nl, loop_DES_rounds_2_xor_31_nl,
          fsm_output(2));
      R_30_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_30_nl, loop_DES_rounds_2_xor_30_nl,
          fsm_output(2));
      R_1_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_29_nl, loop_DES_rounds_2_xor_29_nl,
          fsm_output(2));
      R_29_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_28_nl, loop_DES_rounds_2_xor_28_nl,
          fsm_output(2));
      R_2_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_27_nl, loop_DES_rounds_2_xor_27_nl,
          fsm_output(2));
      R_28_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_26_nl, loop_DES_rounds_2_xor_26_nl,
          fsm_output(2));
      R_3_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_25_nl, loop_DES_rounds_2_xor_25_nl,
          fsm_output(2));
      R_27_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_24_nl, loop_DES_rounds_2_xor_24_nl,
          fsm_output(2));
      R_4_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_23_nl, loop_DES_rounds_2_xor_23_nl,
          fsm_output(2));
      R_26_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_22_nl, loop_DES_rounds_2_xor_22_nl,
          fsm_output(2));
      R_5_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_21_nl, loop_DES_rounds_2_xor_21_nl,
          fsm_output(2));
      R_25_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_20_nl, loop_DES_rounds_2_xor_20_nl,
          fsm_output(2));
      R_6_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_19_nl, loop_DES_rounds_2_xor_19_nl,
          fsm_output(2));
      R_24_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_18_nl, loop_DES_rounds_2_xor_18_nl,
          fsm_output(2));
      R_7_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_17_nl, loop_DES_rounds_2_xor_17_nl,
          fsm_output(2));
      R_23_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_16_nl, loop_DES_rounds_2_xor_16_nl,
          fsm_output(2));
      R_8_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_15_nl, loop_DES_rounds_2_xor_15_nl,
          fsm_output(2));
      R_22_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_14_nl, loop_DES_rounds_2_xor_14_nl,
          fsm_output(2));
      R_9_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_13_nl, loop_DES_rounds_2_xor_13_nl,
          fsm_output(2));
      R_21_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_12_nl, loop_DES_rounds_2_xor_12_nl,
          fsm_output(2));
      R_10_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_11_nl, loop_DES_rounds_2_xor_11_nl,
          fsm_output(2));
      R_20_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_10_nl, loop_DES_rounds_2_xor_10_nl,
          fsm_output(2));
      R_11_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_9_nl, loop_DES_rounds_2_xor_9_nl,
          fsm_output(2));
      R_19_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_8_nl, loop_DES_rounds_2_xor_8_nl,
          fsm_output(2));
      R_12_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_7_nl, loop_DES_rounds_2_xor_7_nl,
          fsm_output(2));
      R_18_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_6_nl, loop_DES_rounds_2_xor_6_nl,
          fsm_output(2));
      R_13_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_5_nl, loop_DES_rounds_2_xor_5_nl,
          fsm_output(2));
      R_17_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_4_nl, loop_DES_rounds_2_xor_4_nl,
          fsm_output(2));
      R_14_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_3_nl, loop_DES_rounds_2_xor_3_nl,
          fsm_output(2));
      R_16_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_2_nl, loop_DES_rounds_2_xor_2_nl,
          fsm_output(2));
      R_15_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_1_nl, loop_DES_rounds_2_xor_1_nl,
          fsm_output(2));
      s_output_1_19_16_5_sva <= operator_8_false_1_read_rom_S_rom_map_1_14_itm;
      s_output_1_3_0_54_sva <= operator_8_false_1_read_rom_S_rom_map_1_13_itm;
      s_output_1_19_16_35_sva <= operator_8_false_1_read_rom_S_rom_map_1_10_itm;
      s_output_1_19_16_20_sva <= operator_8_false_1_read_rom_S_rom_map_1_8_itm;
      s_output_1_3_0_24_sva <= operator_8_false_1_read_rom_S_rom_map_1_9_itm;
      s_output_1_19_16_50_sva <= operator_8_false_1_read_rom_S_rom_map_1_12_itm;
      s_output_1_3_0_39_sva <= operator_8_false_1_read_rom_S_rom_map_1_11_itm;
      s_output_1_3_0_9_sva <= operator_8_false_1_read_rom_S_rom_map_1_15_itm;
      R_24_15_sva <= R_24_13_sva XOR (s_output_1_3_0_37_sva_1(3));
      R_7_15_sva <= R_7_13_sva XOR (s_output_1_3_0_37_sva_1(1));
      R_16_15_sva <= R_16_13_sva XOR (s_output_1_19_16_63_sva_1(2));
      R_15_15_sva <= R_15_13_sva XOR (s_output_1_19_16_33_sva_1(2));
      R_8_15_sva <= R_8_13_sva XOR (s_output_1_19_16_63_sva_1(3));
      R_23_15_sva <= R_23_13_sva XOR (s_output_1_19_16_33_sva_1(3));
      R_0_15_sva <= R_0_13_sva XOR (s_output_1_3_0_67_sva_1(3));
      R_31_15_sva <= R_31_13_sva XOR (s_output_1_19_16_18_sva_1(0));
      R_25_15_sva <= R_25_13_sva XOR (s_output_1_3_0_67_sva_1(0));
      R_6_15_sva <= R_6_13_sva XOR (s_output_1_19_16_18_sva_1(3));
      R_17_15_sva <= R_17_13_sva XOR (s_output_1_3_0_22_sva_1(1));
      R_14_15_sva <= R_14_13_sva XOR (s_output_1_19_16_48_sva_1(0));
      R_9_15_sva <= R_9_13_sva XOR (s_output_1_19_16_33_sva_1(1));
      R_22_15_sva <= R_22_13_sva XOR (s_output_1_19_16_18_sva_1(1));
      R_1_15_sva <= R_1_13_sva XOR (s_output_1_19_16_33_sva_1(0));
      R_30_15_sva <= R_30_13_sva XOR (s_output_1_19_16_48_sva_1(1));
      R_26_15_sva <= R_26_13_sva XOR (s_output_1_19_16_63_sva_1(0));
      R_5_15_sva <= R_5_13_sva XOR (s_output_1_3_0_22_sva_1(2));
      R_18_15_sva <= R_18_13_sva XOR (s_output_1_3_0_37_sva_1(2));
      R_13_15_sva <= R_13_13_sva XOR (s_output_1_3_0_52_sva_1(0));
      R_10_15_sva <= R_10_13_sva XOR (s_output_1_3_0_67_sva_1(1));
      R_21_15_sva <= R_21_13_sva XOR (s_output_1_3_0_52_sva_1(1));
      R_2_15_sva <= R_2_13_sva XOR (s_output_1_19_16_63_sva_1(1));
      R_29_15_sva <= R_29_13_sva XOR (s_output_1_3_0_37_sva_1(0));
      R_27_15_sva <= R_27_13_sva XOR (s_output_1_3_0_22_sva_1(3));
      R_4_15_sva <= R_4_13_sva XOR (s_output_1_19_16_48_sva_1(2));
      R_19_15_sva <= R_19_13_sva XOR (s_output_1_19_16_48_sva_1(3));
      R_12_15_sva <= R_12_13_sva XOR (s_output_1_19_16_18_sva_1(2));
      R_11_15_sva <= R_11_13_sva XOR (s_output_1_3_0_22_sva_1(0));
      R_20_15_sva <= R_20_13_sva XOR (s_output_1_3_0_67_sva_1(2));
      R_3_15_sva <= R_3_13_sva XOR (s_output_1_3_0_52_sva_1(2));
      R_28_15_sva <= R_28_13_sva XOR (s_output_1_3_0_52_sva_1(3));
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_31_3_sva <= R_31_1_sva XOR (s_output_1_19_16_6_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_0_3_sva <= R_0_1_sva XOR (s_output_1_3_0_55_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_30_3_sva <= R_30_1_sva XOR (s_output_1_19_16_36_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_1_3_sva <= R_1_1_sva XOR (s_output_1_19_16_21_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_29_3_sva <= R_29_1_sva XOR (s_output_1_3_0_25_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_2_3_sva <= R_2_1_sva XOR (s_output_1_19_16_51_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_28_3_sva <= R_28_1_sva XOR (s_output_1_3_0_40_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_3_3_sva <= R_3_1_sva XOR (s_output_1_3_0_40_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_27_3_sva <= R_27_1_sva XOR (s_output_1_3_0_10_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_4_3_sva <= R_4_1_sva XOR (s_output_1_19_16_36_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_26_3_sva <= R_26_1_sva XOR (s_output_1_19_16_51_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_5_3_sva <= R_5_1_sva XOR (s_output_1_3_0_10_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_25_3_sva <= R_25_1_sva XOR (s_output_1_3_0_55_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_6_3_sva <= R_6_1_sva XOR (s_output_1_19_16_6_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_24_3_sva <= R_24_1_sva XOR (s_output_1_3_0_25_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_7_3_sva <= R_7_1_sva XOR (s_output_1_3_0_25_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_23_3_sva <= R_23_1_sva XOR (s_output_1_19_16_21_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_8_3_sva <= R_8_1_sva XOR (s_output_1_19_16_51_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_22_3_sva <= R_22_1_sva XOR (s_output_1_19_16_6_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_9_3_sva <= R_9_1_sva XOR (s_output_1_19_16_21_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_21_3_sva <= R_21_1_sva XOR (s_output_1_3_0_40_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_10_3_sva <= R_10_1_sva XOR (s_output_1_3_0_55_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_20_3_sva <= R_20_1_sva XOR (s_output_1_3_0_55_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_11_3_sva <= R_11_1_sva XOR (s_output_1_3_0_10_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_19_3_sva <= R_19_1_sva XOR (s_output_1_19_16_36_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_12_3_sva <= R_12_1_sva XOR (s_output_1_19_16_6_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_18_3_sva <= R_18_1_sva XOR (s_output_1_3_0_25_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_13_3_sva <= R_13_1_sva XOR (s_output_1_3_0_40_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_17_3_sva <= R_17_1_sva XOR (s_output_1_3_0_10_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_14_3_sva <= R_14_1_sva XOR (s_output_1_19_16_36_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_16_3_sva <= R_16_1_sva XOR (s_output_1_19_16_51_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(2)) = '1' ) THEN
        R_15_3_sva <= R_15_1_sva XOR (s_output_1_19_16_21_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_31_4_sva <= R_31_1_sva XOR (s_output_1_19_16_7_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_0_4_sva <= R_0_1_sva XOR (s_output_1_3_0_56_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_30_4_sva <= R_30_1_sva XOR (s_output_1_19_16_37_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_1_4_sva <= R_1_1_sva XOR (s_output_1_19_16_22_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_29_4_sva <= R_29_1_sva XOR (s_output_1_3_0_26_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_2_4_sva <= R_2_1_sva XOR (s_output_1_19_16_52_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_28_4_sva <= R_28_1_sva XOR (s_output_1_3_0_41_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_3_4_sva <= R_3_1_sva XOR (s_output_1_3_0_41_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_27_4_sva <= R_27_1_sva XOR (s_output_1_3_0_11_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_4_4_sva <= R_4_1_sva XOR (s_output_1_19_16_37_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_26_4_sva <= R_26_1_sva XOR (s_output_1_19_16_52_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_5_4_sva <= R_5_1_sva XOR (s_output_1_3_0_11_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_25_4_sva <= R_25_1_sva XOR (s_output_1_3_0_56_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_6_4_sva <= R_6_1_sva XOR (s_output_1_19_16_7_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_24_4_sva <= R_24_1_sva XOR (s_output_1_3_0_26_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_7_4_sva <= R_7_1_sva XOR (s_output_1_3_0_26_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_23_4_sva <= R_23_1_sva XOR (s_output_1_19_16_22_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_8_4_sva <= R_8_1_sva XOR (s_output_1_19_16_52_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_22_4_sva <= R_22_1_sva XOR (s_output_1_19_16_7_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_9_4_sva <= R_9_1_sva XOR (s_output_1_19_16_22_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_21_4_sva <= R_21_1_sva XOR (s_output_1_3_0_41_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_10_4_sva <= R_10_1_sva XOR (s_output_1_3_0_56_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_20_4_sva <= R_20_1_sva XOR (s_output_1_3_0_56_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_11_4_sva <= R_11_1_sva XOR (s_output_1_3_0_11_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_19_4_sva <= R_19_1_sva XOR (s_output_1_19_16_37_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_12_4_sva <= R_12_1_sva XOR (s_output_1_19_16_7_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_18_4_sva <= R_18_1_sva XOR (s_output_1_3_0_26_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_13_4_sva <= R_13_1_sva XOR (s_output_1_3_0_41_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_17_4_sva <= R_17_1_sva XOR (s_output_1_3_0_11_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_14_4_sva <= R_14_1_sva XOR (s_output_1_19_16_37_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_16_4_sva <= R_16_1_sva XOR (s_output_1_19_16_52_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(3)) = '1' ) THEN
        R_15_4_sva <= R_15_1_sva XOR (s_output_1_19_16_22_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_31_5_sva <= R_31_3_sva XOR (s_output_1_19_16_8_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_0_5_sva <= R_0_3_sva XOR (s_output_1_3_0_57_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_30_5_sva <= R_30_3_sva XOR (s_output_1_19_16_38_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_1_5_sva <= R_1_3_sva XOR (s_output_1_19_16_23_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_29_5_sva <= R_29_3_sva XOR (s_output_1_3_0_27_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_2_5_sva <= R_2_3_sva XOR (s_output_1_19_16_53_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_28_5_sva <= R_28_3_sva XOR (s_output_1_3_0_42_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_3_5_sva <= R_3_3_sva XOR (s_output_1_3_0_42_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_27_5_sva <= R_27_3_sva XOR (s_output_1_3_0_12_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_4_5_sva <= R_4_3_sva XOR (s_output_1_19_16_38_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_26_5_sva <= R_26_3_sva XOR (s_output_1_19_16_53_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_5_5_sva <= R_5_3_sva XOR (s_output_1_3_0_12_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_25_5_sva <= R_25_3_sva XOR (s_output_1_3_0_57_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_6_5_sva <= R_6_3_sva XOR (s_output_1_19_16_8_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_24_5_sva <= R_24_3_sva XOR (s_output_1_3_0_27_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_7_5_sva <= R_7_3_sva XOR (s_output_1_3_0_27_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_23_5_sva <= R_23_3_sva XOR (s_output_1_19_16_23_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_8_5_sva <= R_8_3_sva XOR (s_output_1_19_16_53_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_22_5_sva <= R_22_3_sva XOR (s_output_1_19_16_8_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_9_5_sva <= R_9_3_sva XOR (s_output_1_19_16_23_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_21_5_sva <= R_21_3_sva XOR (s_output_1_3_0_42_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_10_5_sva <= R_10_3_sva XOR (s_output_1_3_0_57_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_20_5_sva <= R_20_3_sva XOR (s_output_1_3_0_57_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_11_5_sva <= R_11_3_sva XOR (s_output_1_3_0_12_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_19_5_sva <= R_19_3_sva XOR (s_output_1_19_16_38_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_12_5_sva <= R_12_3_sva XOR (s_output_1_19_16_8_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_18_5_sva <= R_18_3_sva XOR (s_output_1_3_0_27_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_13_5_sva <= R_13_3_sva XOR (s_output_1_3_0_42_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_17_5_sva <= R_17_3_sva XOR (s_output_1_3_0_12_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_14_5_sva <= R_14_3_sva XOR (s_output_1_19_16_38_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_16_5_sva <= R_16_3_sva XOR (s_output_1_19_16_53_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '1' ) THEN
        R_15_5_sva <= R_15_3_sva XOR (s_output_1_19_16_23_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_31_6_sva <= R_31_4_sva XOR (s_output_1_19_16_9_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_0_6_sva <= R_0_4_sva XOR (s_output_1_3_0_58_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_30_6_sva <= R_30_4_sva XOR (s_output_1_19_16_39_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_1_6_sva <= R_1_4_sva XOR (s_output_1_19_16_24_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_29_6_sva <= R_29_4_sva XOR (s_output_1_3_0_28_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_2_6_sva <= R_2_4_sva XOR (s_output_1_19_16_54_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_28_6_sva <= R_28_4_sva XOR (s_output_1_3_0_43_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_3_6_sva <= R_3_4_sva XOR (s_output_1_3_0_43_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_27_6_sva <= R_27_4_sva XOR (s_output_1_3_0_13_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_4_6_sva <= R_4_4_sva XOR (s_output_1_19_16_39_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_26_6_sva <= R_26_4_sva XOR (s_output_1_19_16_54_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_5_6_sva <= R_5_4_sva XOR (s_output_1_3_0_13_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_25_6_sva <= R_25_4_sva XOR (s_output_1_3_0_58_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_6_6_sva <= R_6_4_sva XOR (s_output_1_19_16_9_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_24_6_sva <= R_24_4_sva XOR (s_output_1_3_0_28_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_7_6_sva <= R_7_4_sva XOR (s_output_1_3_0_28_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_23_6_sva <= R_23_4_sva XOR (s_output_1_19_16_24_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_8_6_sva <= R_8_4_sva XOR (s_output_1_19_16_54_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_22_6_sva <= R_22_4_sva XOR (s_output_1_19_16_9_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_9_6_sva <= R_9_4_sva XOR (s_output_1_19_16_24_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_21_6_sva <= R_21_4_sva XOR (s_output_1_3_0_43_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_10_6_sva <= R_10_4_sva XOR (s_output_1_3_0_58_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_20_6_sva <= R_20_4_sva XOR (s_output_1_3_0_58_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_11_6_sva <= R_11_4_sva XOR (s_output_1_3_0_13_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_19_6_sva <= R_19_4_sva XOR (s_output_1_19_16_39_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_12_6_sva <= R_12_4_sva XOR (s_output_1_19_16_9_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_18_6_sva <= R_18_4_sva XOR (s_output_1_3_0_28_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_13_6_sva <= R_13_4_sva XOR (s_output_1_3_0_43_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_17_6_sva <= R_17_4_sva XOR (s_output_1_3_0_13_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_14_6_sva <= R_14_4_sva XOR (s_output_1_19_16_39_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_16_6_sva <= R_16_4_sva XOR (s_output_1_19_16_54_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(5)) = '1' ) THEN
        R_15_6_sva <= R_15_4_sva XOR (s_output_1_19_16_24_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_31_7_sva <= R_31_5_sva XOR (s_output_1_19_16_10_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_0_7_sva <= R_0_5_sva XOR (s_output_1_3_0_59_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_30_7_sva <= R_30_5_sva XOR (s_output_1_19_16_40_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_1_7_sva <= R_1_5_sva XOR (s_output_1_19_16_25_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_29_7_sva <= R_29_5_sva XOR (s_output_1_3_0_29_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_2_7_sva <= R_2_5_sva XOR (s_output_1_19_16_55_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_28_7_sva <= R_28_5_sva XOR (s_output_1_3_0_44_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_3_7_sva <= R_3_5_sva XOR (s_output_1_3_0_44_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_27_7_sva <= R_27_5_sva XOR (s_output_1_3_0_14_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_4_7_sva <= R_4_5_sva XOR (s_output_1_19_16_40_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_26_7_sva <= R_26_5_sva XOR (s_output_1_19_16_55_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_5_7_sva <= R_5_5_sva XOR (s_output_1_3_0_14_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_25_7_sva <= R_25_5_sva XOR (s_output_1_3_0_59_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_6_7_sva <= R_6_5_sva XOR (s_output_1_19_16_10_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_24_7_sva <= R_24_5_sva XOR (s_output_1_3_0_29_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_7_7_sva <= R_7_5_sva XOR (s_output_1_3_0_29_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_23_7_sva <= R_23_5_sva XOR (s_output_1_19_16_25_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_8_7_sva <= R_8_5_sva XOR (s_output_1_19_16_55_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_22_7_sva <= R_22_5_sva XOR (s_output_1_19_16_10_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_9_7_sva <= R_9_5_sva XOR (s_output_1_19_16_25_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_21_7_sva <= R_21_5_sva XOR (s_output_1_3_0_44_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_10_7_sva <= R_10_5_sva XOR (s_output_1_3_0_59_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_20_7_sva <= R_20_5_sva XOR (s_output_1_3_0_59_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_11_7_sva <= R_11_5_sva XOR (s_output_1_3_0_14_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_19_7_sva <= R_19_5_sva XOR (s_output_1_19_16_40_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_12_7_sva <= R_12_5_sva XOR (s_output_1_19_16_10_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_18_7_sva <= R_18_5_sva XOR (s_output_1_3_0_29_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_13_7_sva <= R_13_5_sva XOR (s_output_1_3_0_44_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_17_7_sva <= R_17_5_sva XOR (s_output_1_3_0_14_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_14_7_sva <= R_14_5_sva XOR (s_output_1_19_16_40_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_16_7_sva <= R_16_5_sva XOR (s_output_1_19_16_55_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(6)) = '1' ) THEN
        R_15_7_sva <= R_15_5_sva XOR (s_output_1_19_16_25_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_31_8_sva <= R_31_6_sva XOR (s_output_1_19_16_11_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_0_8_sva <= R_0_6_sva XOR (s_output_1_3_0_60_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_30_8_sva <= R_30_6_sva XOR (s_output_1_19_16_41_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_1_8_sva <= R_1_6_sva XOR (s_output_1_19_16_26_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_29_8_sva <= R_29_6_sva XOR (s_output_1_3_0_30_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_2_8_sva <= R_2_6_sva XOR (s_output_1_19_16_56_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_28_8_sva <= R_28_6_sva XOR (s_output_1_3_0_45_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_3_8_sva <= R_3_6_sva XOR (s_output_1_3_0_45_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_27_8_sva <= R_27_6_sva XOR (s_output_1_3_0_15_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_4_8_sva <= R_4_6_sva XOR (s_output_1_19_16_41_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_26_8_sva <= R_26_6_sva XOR (s_output_1_19_16_56_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_5_8_sva <= R_5_6_sva XOR (s_output_1_3_0_15_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_25_8_sva <= R_25_6_sva XOR (s_output_1_3_0_60_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_6_8_sva <= R_6_6_sva XOR (s_output_1_19_16_11_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_24_8_sva <= R_24_6_sva XOR (s_output_1_3_0_30_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_7_8_sva <= R_7_6_sva XOR (s_output_1_3_0_30_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_23_8_sva <= R_23_6_sva XOR (s_output_1_19_16_26_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_8_8_sva <= R_8_6_sva XOR (s_output_1_19_16_56_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_22_8_sva <= R_22_6_sva XOR (s_output_1_19_16_11_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_9_8_sva <= R_9_6_sva XOR (s_output_1_19_16_26_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_21_8_sva <= R_21_6_sva XOR (s_output_1_3_0_45_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_10_8_sva <= R_10_6_sva XOR (s_output_1_3_0_60_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_20_8_sva <= R_20_6_sva XOR (s_output_1_3_0_60_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_11_8_sva <= R_11_6_sva XOR (s_output_1_3_0_15_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_19_8_sva <= R_19_6_sva XOR (s_output_1_19_16_41_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_12_8_sva <= R_12_6_sva XOR (s_output_1_19_16_11_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_18_8_sva <= R_18_6_sva XOR (s_output_1_3_0_30_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_13_8_sva <= R_13_6_sva XOR (s_output_1_3_0_45_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_17_8_sva <= R_17_6_sva XOR (s_output_1_3_0_15_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_14_8_sva <= R_14_6_sva XOR (s_output_1_19_16_41_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_16_8_sva <= R_16_6_sva XOR (s_output_1_19_16_56_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(7)) = '1' ) THEN
        R_15_8_sva <= R_15_6_sva XOR (s_output_1_19_16_26_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_31_9_sva <= R_31_7_sva XOR (s_output_1_19_16_12_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_0_9_sva <= R_0_7_sva XOR (s_output_1_3_0_61_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_30_9_sva <= R_30_7_sva XOR (s_output_1_19_16_42_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_1_9_sva <= R_1_7_sva XOR (s_output_1_19_16_27_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_29_9_sva <= R_29_7_sva XOR (s_output_1_3_0_31_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_2_9_sva <= R_2_7_sva XOR (s_output_1_19_16_57_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_28_9_sva <= R_28_7_sva XOR (s_output_1_3_0_46_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_3_9_sva <= R_3_7_sva XOR (s_output_1_3_0_46_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_27_9_sva <= R_27_7_sva XOR (s_output_1_3_0_16_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_4_9_sva <= R_4_7_sva XOR (s_output_1_19_16_42_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_26_9_sva <= R_26_7_sva XOR (s_output_1_19_16_57_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_5_9_sva <= R_5_7_sva XOR (s_output_1_3_0_16_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_25_9_sva <= R_25_7_sva XOR (s_output_1_3_0_61_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_6_9_sva <= R_6_7_sva XOR (s_output_1_19_16_12_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_24_9_sva <= R_24_7_sva XOR (s_output_1_3_0_31_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_7_9_sva <= R_7_7_sva XOR (s_output_1_3_0_31_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_23_9_sva <= R_23_7_sva XOR (s_output_1_19_16_27_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_8_9_sva <= R_8_7_sva XOR (s_output_1_19_16_57_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_22_9_sva <= R_22_7_sva XOR (s_output_1_19_16_12_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_9_9_sva <= R_9_7_sva XOR (s_output_1_19_16_27_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_21_9_sva <= R_21_7_sva XOR (s_output_1_3_0_46_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_10_9_sva <= R_10_7_sva XOR (s_output_1_3_0_61_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_20_9_sva <= R_20_7_sva XOR (s_output_1_3_0_61_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_11_9_sva <= R_11_7_sva XOR (s_output_1_3_0_16_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_19_9_sva <= R_19_7_sva XOR (s_output_1_19_16_42_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_12_9_sva <= R_12_7_sva XOR (s_output_1_19_16_12_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_18_9_sva <= R_18_7_sva XOR (s_output_1_3_0_31_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_13_9_sva <= R_13_7_sva XOR (s_output_1_3_0_46_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_17_9_sva <= R_17_7_sva XOR (s_output_1_3_0_16_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_14_9_sva <= R_14_7_sva XOR (s_output_1_19_16_42_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_16_9_sva <= R_16_7_sva XOR (s_output_1_19_16_57_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(8)) = '1' ) THEN
        R_15_9_sva <= R_15_7_sva XOR (s_output_1_19_16_27_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_31_10_sva <= R_31_8_sva XOR (s_output_1_19_16_13_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_0_10_sva <= R_0_8_sva XOR (s_output_1_3_0_62_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_30_10_sva <= R_30_8_sva XOR (s_output_1_19_16_43_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_1_10_sva <= R_1_8_sva XOR (s_output_1_19_16_28_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_29_10_sva <= R_29_8_sva XOR (s_output_1_3_0_32_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_2_10_sva <= R_2_8_sva XOR (s_output_1_19_16_58_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_28_10_sva <= R_28_8_sva XOR (s_output_1_3_0_47_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_3_10_sva <= R_3_8_sva XOR (s_output_1_3_0_47_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_27_10_sva <= R_27_8_sva XOR (s_output_1_3_0_17_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_4_10_sva <= R_4_8_sva XOR (s_output_1_19_16_43_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_26_10_sva <= R_26_8_sva XOR (s_output_1_19_16_58_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_5_10_sva <= R_5_8_sva XOR (s_output_1_3_0_17_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_25_10_sva <= R_25_8_sva XOR (s_output_1_3_0_62_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_6_10_sva <= R_6_8_sva XOR (s_output_1_19_16_13_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_24_10_sva <= R_24_8_sva XOR (s_output_1_3_0_32_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_7_10_sva <= R_7_8_sva XOR (s_output_1_3_0_32_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_23_10_sva <= R_23_8_sva XOR (s_output_1_19_16_28_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_8_10_sva <= R_8_8_sva XOR (s_output_1_19_16_58_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_22_10_sva <= R_22_8_sva XOR (s_output_1_19_16_13_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_9_10_sva <= R_9_8_sva XOR (s_output_1_19_16_28_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_21_10_sva <= R_21_8_sva XOR (s_output_1_3_0_47_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_10_10_sva <= R_10_8_sva XOR (s_output_1_3_0_62_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_20_10_sva <= R_20_8_sva XOR (s_output_1_3_0_62_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_11_10_sva <= R_11_8_sva XOR (s_output_1_3_0_17_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_19_10_sva <= R_19_8_sva XOR (s_output_1_19_16_43_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_12_10_sva <= R_12_8_sva XOR (s_output_1_19_16_13_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_18_10_sva <= R_18_8_sva XOR (s_output_1_3_0_32_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_13_10_sva <= R_13_8_sva XOR (s_output_1_3_0_47_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_17_10_sva <= R_17_8_sva XOR (s_output_1_3_0_17_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_14_10_sva <= R_14_8_sva XOR (s_output_1_19_16_43_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_16_10_sva <= R_16_8_sva XOR (s_output_1_19_16_58_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(9)) = '1' ) THEN
        R_15_10_sva <= R_15_8_sva XOR (s_output_1_19_16_28_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_31_11_sva <= R_31_9_sva XOR (s_output_1_19_16_14_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_0_11_sva <= R_0_9_sva XOR (s_output_1_3_0_63_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_30_11_sva <= R_30_9_sva XOR (s_output_1_19_16_44_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_1_11_sva <= R_1_9_sva XOR (s_output_1_19_16_29_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_29_11_sva <= R_29_9_sva XOR (s_output_1_3_0_33_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_2_11_sva <= R_2_9_sva XOR (s_output_1_19_16_59_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_28_11_sva <= R_28_9_sva XOR (s_output_1_3_0_48_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_3_11_sva <= R_3_9_sva XOR (s_output_1_3_0_48_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_27_11_sva <= R_27_9_sva XOR (s_output_1_3_0_18_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_4_11_sva <= R_4_9_sva XOR (s_output_1_19_16_44_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_26_11_sva <= R_26_9_sva XOR (s_output_1_19_16_59_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_5_11_sva <= R_5_9_sva XOR (s_output_1_3_0_18_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_25_11_sva <= R_25_9_sva XOR (s_output_1_3_0_63_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_6_11_sva <= R_6_9_sva XOR (s_output_1_19_16_14_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_24_11_sva <= R_24_9_sva XOR (s_output_1_3_0_33_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_7_11_sva <= R_7_9_sva XOR (s_output_1_3_0_33_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_23_11_sva <= R_23_9_sva XOR (s_output_1_19_16_29_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_8_11_sva <= R_8_9_sva XOR (s_output_1_19_16_59_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_22_11_sva <= R_22_9_sva XOR (s_output_1_19_16_14_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_9_11_sva <= R_9_9_sva XOR (s_output_1_19_16_29_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_21_11_sva <= R_21_9_sva XOR (s_output_1_3_0_48_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_10_11_sva <= R_10_9_sva XOR (s_output_1_3_0_63_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_20_11_sva <= R_20_9_sva XOR (s_output_1_3_0_63_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_11_11_sva <= R_11_9_sva XOR (s_output_1_3_0_18_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_19_11_sva <= R_19_9_sva XOR (s_output_1_19_16_44_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_12_11_sva <= R_12_9_sva XOR (s_output_1_19_16_14_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_18_11_sva <= R_18_9_sva XOR (s_output_1_3_0_33_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_13_11_sva <= R_13_9_sva XOR (s_output_1_3_0_48_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_17_11_sva <= R_17_9_sva XOR (s_output_1_3_0_18_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_14_11_sva <= R_14_9_sva XOR (s_output_1_19_16_44_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_16_11_sva <= R_16_9_sva XOR (s_output_1_19_16_59_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(10)) = '1' ) THEN
        R_15_11_sva <= R_15_9_sva XOR (s_output_1_19_16_29_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_31_12_sva <= R_31_10_sva XOR (s_output_1_19_16_15_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_0_12_sva <= R_0_10_sva XOR (s_output_1_3_0_64_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_30_12_sva <= R_30_10_sva XOR (s_output_1_19_16_45_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_1_12_sva <= R_1_10_sva XOR (s_output_1_19_16_30_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_29_12_sva <= R_29_10_sva XOR (s_output_1_3_0_34_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_2_12_sva <= R_2_10_sva XOR (s_output_1_19_16_60_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_28_12_sva <= R_28_10_sva XOR (s_output_1_3_0_49_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_3_12_sva <= R_3_10_sva XOR (s_output_1_3_0_49_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_27_12_sva <= R_27_10_sva XOR (s_output_1_3_0_19_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_4_12_sva <= R_4_10_sva XOR (s_output_1_19_16_45_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_26_12_sva <= R_26_10_sva XOR (s_output_1_19_16_60_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_5_12_sva <= R_5_10_sva XOR (s_output_1_3_0_19_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_25_12_sva <= R_25_10_sva XOR (s_output_1_3_0_64_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_6_12_sva <= R_6_10_sva XOR (s_output_1_19_16_15_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_24_12_sva <= R_24_10_sva XOR (s_output_1_3_0_34_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_7_12_sva <= R_7_10_sva XOR (s_output_1_3_0_34_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_23_12_sva <= R_23_10_sva XOR (s_output_1_19_16_30_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_8_12_sva <= R_8_10_sva XOR (s_output_1_19_16_60_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_22_12_sva <= R_22_10_sva XOR (s_output_1_19_16_15_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_9_12_sva <= R_9_10_sva XOR (s_output_1_19_16_30_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_21_12_sva <= R_21_10_sva XOR (s_output_1_3_0_49_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_10_12_sva <= R_10_10_sva XOR (s_output_1_3_0_64_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_20_12_sva <= R_20_10_sva XOR (s_output_1_3_0_64_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_11_12_sva <= R_11_10_sva XOR (s_output_1_3_0_19_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_19_12_sva <= R_19_10_sva XOR (s_output_1_19_16_45_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_12_12_sva <= R_12_10_sva XOR (s_output_1_19_16_15_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_18_12_sva <= R_18_10_sva XOR (s_output_1_3_0_34_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_13_12_sva <= R_13_10_sva XOR (s_output_1_3_0_49_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_17_12_sva <= R_17_10_sva XOR (s_output_1_3_0_19_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_14_12_sva <= R_14_10_sva XOR (s_output_1_19_16_45_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_16_12_sva <= R_16_10_sva XOR (s_output_1_19_16_60_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(11)) = '1' ) THEN
        R_15_12_sva <= R_15_10_sva XOR (s_output_1_19_16_30_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_31_13_sva <= R_31_11_sva XOR (s_output_1_19_16_16_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_0_13_sva <= R_0_11_sva XOR (s_output_1_3_0_65_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_30_13_sva <= R_30_11_sva XOR (s_output_1_19_16_46_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_1_13_sva <= R_1_11_sva XOR (s_output_1_19_16_31_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_29_13_sva <= R_29_11_sva XOR (s_output_1_3_0_35_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_2_13_sva <= R_2_11_sva XOR (s_output_1_19_16_61_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_28_13_sva <= R_28_11_sva XOR (s_output_1_3_0_50_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_3_13_sva <= R_3_11_sva XOR (s_output_1_3_0_50_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_27_13_sva <= R_27_11_sva XOR (s_output_1_3_0_20_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_4_13_sva <= R_4_11_sva XOR (s_output_1_19_16_46_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_26_13_sva <= R_26_11_sva XOR (s_output_1_19_16_61_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_5_13_sva <= R_5_11_sva XOR (s_output_1_3_0_20_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_25_13_sva <= R_25_11_sva XOR (s_output_1_3_0_65_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_6_13_sva <= R_6_11_sva XOR (s_output_1_19_16_16_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_24_13_sva <= R_24_11_sva XOR (s_output_1_3_0_35_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_7_13_sva <= R_7_11_sva XOR (s_output_1_3_0_35_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_23_13_sva <= R_23_11_sva XOR (s_output_1_19_16_31_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_8_13_sva <= R_8_11_sva XOR (s_output_1_19_16_61_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_22_13_sva <= R_22_11_sva XOR (s_output_1_19_16_16_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_9_13_sva <= R_9_11_sva XOR (s_output_1_19_16_31_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_21_13_sva <= R_21_11_sva XOR (s_output_1_3_0_50_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_10_13_sva <= R_10_11_sva XOR (s_output_1_3_0_65_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_20_13_sva <= R_20_11_sva XOR (s_output_1_3_0_65_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_11_13_sva <= R_11_11_sva XOR (s_output_1_3_0_20_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_19_13_sva <= R_19_11_sva XOR (s_output_1_19_16_46_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_12_13_sva <= R_12_11_sva XOR (s_output_1_19_16_16_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_18_13_sva <= R_18_11_sva XOR (s_output_1_3_0_35_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_13_13_sva <= R_13_11_sva XOR (s_output_1_3_0_50_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_17_13_sva <= R_17_11_sva XOR (s_output_1_3_0_20_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_14_13_sva <= R_14_11_sva XOR (s_output_1_19_16_46_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_16_13_sva <= R_16_11_sva XOR (s_output_1_19_16_61_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(12)) = '1' ) THEN
        R_15_13_sva <= R_15_11_sva XOR (s_output_1_19_16_31_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_7_14_sva <= R_7_12_sva XOR (s_output_1_3_0_36_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_24_14_sva <= R_24_12_sva XOR (s_output_1_3_0_36_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_15_14_sva <= R_15_12_sva XOR (s_output_1_19_16_32_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_16_14_sva <= R_16_12_sva XOR (s_output_1_19_16_62_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_23_14_sva <= R_23_12_sva XOR (s_output_1_19_16_32_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_8_14_sva <= R_8_12_sva XOR (s_output_1_19_16_62_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_31_14_sva <= R_31_12_sva XOR (s_output_1_19_16_17_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_0_14_sva <= R_0_12_sva XOR (s_output_1_3_0_66_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_6_14_sva <= R_6_12_sva XOR (s_output_1_19_16_17_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_25_14_sva <= R_25_12_sva XOR (s_output_1_3_0_66_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_14_14_sva <= R_14_12_sva XOR (s_output_1_19_16_47_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_17_14_sva <= R_17_12_sva XOR (s_output_1_3_0_21_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_22_14_sva <= R_22_12_sva XOR (s_output_1_19_16_17_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_9_14_sva <= R_9_12_sva XOR (s_output_1_19_16_32_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_30_14_sva <= R_30_12_sva XOR (s_output_1_19_16_47_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_1_14_sva <= R_1_12_sva XOR (s_output_1_19_16_32_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_5_14_sva <= R_5_12_sva XOR (s_output_1_3_0_21_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_26_14_sva <= R_26_12_sva XOR (s_output_1_19_16_62_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_13_14_sva <= R_13_12_sva XOR (s_output_1_3_0_51_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_18_14_sva <= R_18_12_sva XOR (s_output_1_3_0_36_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_21_14_sva <= R_21_12_sva XOR (s_output_1_3_0_51_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_10_14_sva <= R_10_12_sva XOR (s_output_1_3_0_66_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_29_14_sva <= R_29_12_sva XOR (s_output_1_3_0_36_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_2_14_sva <= R_2_12_sva XOR (s_output_1_19_16_62_sva_1(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_4_14_sva <= R_4_12_sva XOR (s_output_1_19_16_47_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_27_14_sva <= R_27_12_sva XOR (s_output_1_3_0_21_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_12_14_sva <= R_12_12_sva XOR (s_output_1_19_16_17_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_19_14_sva <= R_19_12_sva XOR (s_output_1_19_16_47_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_20_14_sva <= R_20_12_sva XOR (s_output_1_3_0_66_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_11_14_sva <= R_11_12_sva XOR (s_output_1_3_0_21_sva_1(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_28_14_sva <= R_28_12_sva XOR (s_output_1_3_0_51_sva_1(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(13)) = '1' ) THEN
        R_3_14_sva <= R_3_12_sva XOR (s_output_1_3_0_51_sva_1(2));
      END IF;
    END IF;
  END PROCESS;
  loop_DES_rounds_1_xor_32_nl <= (input_sva(6)) XOR (s_output_1_19_16_4_sva(0));
  loop_DES_rounds_2_xor_32_nl <= (input_sva(7)) XOR (s_output_1_19_16_5_sva(0));
  loop_DES_rounds_1_xor_31_nl <= (input_sva(56)) XOR (s_output_1_3_0_53_sva(3));
  loop_DES_rounds_2_xor_31_nl <= (input_sva(57)) XOR (s_output_1_3_0_54_sva(3));
  loop_DES_rounds_1_xor_30_nl <= (input_sva(14)) XOR (s_output_1_19_16_34_sva(1));
  loop_DES_rounds_2_xor_30_nl <= (input_sva(15)) XOR (s_output_1_19_16_35_sva(1));
  loop_DES_rounds_1_xor_29_nl <= (input_sva(48)) XOR (s_output_1_19_16_19_sva(0));
  loop_DES_rounds_2_xor_29_nl <= (input_sva(49)) XOR (s_output_1_19_16_20_sva(0));
  loop_DES_rounds_1_xor_28_nl <= (input_sva(22)) XOR (s_output_1_3_0_23_sva(0));
  loop_DES_rounds_2_xor_28_nl <= (input_sva(23)) XOR (s_output_1_3_0_24_sva(0));
  loop_DES_rounds_1_xor_27_nl <= (input_sva(40)) XOR (s_output_1_19_16_49_sva(1));
  loop_DES_rounds_2_xor_27_nl <= (input_sva(41)) XOR (s_output_1_19_16_50_sva(1));
  loop_DES_rounds_1_xor_26_nl <= (input_sva(30)) XOR (s_output_1_3_0_38_sva(3));
  loop_DES_rounds_2_xor_26_nl <= (input_sva(31)) XOR (s_output_1_3_0_39_sva(3));
  loop_DES_rounds_1_xor_25_nl <= (input_sva(32)) XOR (s_output_1_3_0_38_sva(2));
  loop_DES_rounds_2_xor_25_nl <= (input_sva(33)) XOR (s_output_1_3_0_39_sva(2));
  loop_DES_rounds_1_xor_24_nl <= (input_sva(38)) XOR (s_output_1_3_0_8_sva(3));
  loop_DES_rounds_2_xor_24_nl <= (input_sva(39)) XOR (s_output_1_3_0_9_sva(3));
  loop_DES_rounds_1_xor_23_nl <= (input_sva(24)) XOR (s_output_1_19_16_34_sva(2));
  loop_DES_rounds_2_xor_23_nl <= (input_sva(25)) XOR (s_output_1_19_16_35_sva(2));
  loop_DES_rounds_1_xor_22_nl <= (input_sva(46)) XOR (s_output_1_19_16_49_sva(0));
  loop_DES_rounds_2_xor_22_nl <= (input_sva(47)) XOR (s_output_1_19_16_50_sva(0));
  loop_DES_rounds_1_xor_21_nl <= (input_sva(16)) XOR (s_output_1_3_0_8_sva(2));
  loop_DES_rounds_2_xor_21_nl <= (input_sva(17)) XOR (s_output_1_3_0_9_sva(2));
  loop_DES_rounds_1_xor_20_nl <= (input_sva(54)) XOR (s_output_1_3_0_53_sva(0));
  loop_DES_rounds_2_xor_20_nl <= (input_sva(55)) XOR (s_output_1_3_0_54_sva(0));
  loop_DES_rounds_1_xor_19_nl <= (input_sva(8)) XOR (s_output_1_19_16_4_sva(3));
  loop_DES_rounds_2_xor_19_nl <= (input_sva(9)) XOR (s_output_1_19_16_5_sva(3));
  loop_DES_rounds_1_xor_18_nl <= (input_sva(62)) XOR (s_output_1_3_0_23_sva(3));
  loop_DES_rounds_2_xor_18_nl <= (input_sva(63)) XOR (s_output_1_3_0_24_sva(3));
  loop_DES_rounds_1_xor_17_nl <= (input_sva(0)) XOR (s_output_1_3_0_23_sva(1));
  loop_DES_rounds_2_xor_17_nl <= (input_sva(1)) XOR (s_output_1_3_0_24_sva(1));
  loop_DES_rounds_1_xor_16_nl <= (input_sva(4)) XOR (s_output_1_19_16_19_sva(3));
  loop_DES_rounds_2_xor_16_nl <= (input_sva(5)) XOR (s_output_1_19_16_20_sva(3));
  loop_DES_rounds_1_xor_15_nl <= (input_sva(58)) XOR (s_output_1_19_16_49_sva(3));
  loop_DES_rounds_2_xor_15_nl <= (input_sva(59)) XOR (s_output_1_19_16_50_sva(3));
  loop_DES_rounds_1_xor_14_nl <= (input_sva(12)) XOR (s_output_1_19_16_4_sva(1));
  loop_DES_rounds_2_xor_14_nl <= (input_sva(13)) XOR (s_output_1_19_16_5_sva(1));
  loop_DES_rounds_1_xor_13_nl <= (input_sva(50)) XOR (s_output_1_19_16_19_sva(1));
  loop_DES_rounds_2_xor_13_nl <= (input_sva(51)) XOR (s_output_1_19_16_20_sva(1));
  loop_DES_rounds_1_xor_12_nl <= (input_sva(20)) XOR (s_output_1_3_0_38_sva(1));
  loop_DES_rounds_2_xor_12_nl <= (input_sva(21)) XOR (s_output_1_3_0_39_sva(1));
  loop_DES_rounds_1_xor_11_nl <= (input_sva(42)) XOR (s_output_1_3_0_53_sva(1));
  loop_DES_rounds_2_xor_11_nl <= (input_sva(43)) XOR (s_output_1_3_0_54_sva(1));
  loop_DES_rounds_1_xor_10_nl <= (input_sva(28)) XOR (s_output_1_3_0_53_sva(2));
  loop_DES_rounds_2_xor_10_nl <= (input_sva(29)) XOR (s_output_1_3_0_54_sva(2));
  loop_DES_rounds_1_xor_9_nl <= (input_sva(34)) XOR (s_output_1_3_0_8_sva(0));
  loop_DES_rounds_2_xor_9_nl <= (input_sva(35)) XOR (s_output_1_3_0_9_sva(0));
  loop_DES_rounds_1_xor_8_nl <= (input_sva(36)) XOR (s_output_1_19_16_34_sva(3));
  loop_DES_rounds_2_xor_8_nl <= (input_sva(37)) XOR (s_output_1_19_16_35_sva(3));
  loop_DES_rounds_1_xor_7_nl <= (input_sva(26)) XOR (s_output_1_19_16_4_sva(2));
  loop_DES_rounds_2_xor_7_nl <= (input_sva(27)) XOR (s_output_1_19_16_5_sva(2));
  loop_DES_rounds_1_xor_6_nl <= (input_sva(44)) XOR (s_output_1_3_0_23_sva(2));
  loop_DES_rounds_2_xor_6_nl <= (input_sva(45)) XOR (s_output_1_3_0_24_sva(2));
  loop_DES_rounds_1_xor_5_nl <= (input_sva(18)) XOR (s_output_1_3_0_38_sva(0));
  loop_DES_rounds_2_xor_5_nl <= (input_sva(19)) XOR (s_output_1_3_0_39_sva(0));
  loop_DES_rounds_1_xor_4_nl <= (input_sva(52)) XOR (s_output_1_3_0_8_sva(1));
  loop_DES_rounds_2_xor_4_nl <= (input_sva(53)) XOR (s_output_1_3_0_9_sva(1));
  loop_DES_rounds_1_xor_3_nl <= (input_sva(10)) XOR (s_output_1_19_16_34_sva(0));
  loop_DES_rounds_2_xor_3_nl <= (input_sva(11)) XOR (s_output_1_19_16_35_sva(0));
  loop_DES_rounds_1_xor_2_nl <= (input_sva(60)) XOR (s_output_1_19_16_49_sva(2));
  loop_DES_rounds_2_xor_2_nl <= (input_sva(61)) XOR (s_output_1_19_16_50_sva(2));
  loop_DES_rounds_1_xor_1_nl <= (input_sva(2)) XOR (s_output_1_19_16_19_sva(2));
  loop_DES_rounds_2_xor_1_nl <= (input_sva(3)) XOR (s_output_1_19_16_20_sva(2));
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    des_check
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;


ENTITY des_check IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    input_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    input_rsc_triosy_lz : OUT STD_LOGIC;
    key_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    key_rsc_triosy_lz : OUT STD_LOGIC;
    return_rsc_dat : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    return_rsc_triosy_lz : OUT STD_LOGIC
  );
END des_check;

ARCHITECTURE v1 OF des_check IS
  -- Default Constants

  COMPONENT des_check_core
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      input_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      input_rsc_triosy_lz : OUT STD_LOGIC;
      key_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      key_rsc_triosy_lz : OUT STD_LOGIC;
      return_rsc_dat : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      return_rsc_triosy_lz : OUT STD_LOGIC
    );
  END COMPONENT;
  SIGNAL des_check_core_inst_input_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL des_check_core_inst_key_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL des_check_core_inst_return_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  des_check_core_inst : des_check_core
    PORT MAP(
      clk => clk,
      rst => rst,
      input_rsc_dat => des_check_core_inst_input_rsc_dat,
      input_rsc_triosy_lz => input_rsc_triosy_lz,
      key_rsc_dat => des_check_core_inst_key_rsc_dat,
      key_rsc_triosy_lz => key_rsc_triosy_lz,
      return_rsc_dat => des_check_core_inst_return_rsc_dat,
      return_rsc_triosy_lz => return_rsc_triosy_lz
    );
  des_check_core_inst_input_rsc_dat <= input_rsc_dat;
  des_check_core_inst_key_rsc_dat <= key_rsc_dat;
  return_rsc_dat <= des_check_core_inst_return_rsc_dat;

END v1;



