
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl_des_checkmgc_rom_12_512_4_1.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Sun Mar 21 12:44:05 2021
// ----------------------------------------------------------------------

// 
module des_checkmgc_rom_12_512_4_1 (addr, data_out
);
  input [8:0]addr ;
  output [3:0]data_out ;


  // Constants for ROM dimensions
  parameter n_width    = 4;
  parameter n_size     = 512;
  parameter n_numports = 1;
  parameter n_addr_w   = 9;
  parameter n_inreg    = 0;
  parameter n_outreg   = 0;

  // Declare storage for memory elements
  (* rom_style = "block" *)
  wire [3:0] mem [511:0];

  // Declare output registers
  reg [3:0] data_out_t;

  // Initialize ROM contents
  // pragma attribute mem rom_block TRUE
  assign mem[0] = 4'b1110;
  assign mem[1] = 4'b0100;
  assign mem[2] = 4'b1101;
  assign mem[3] = 4'b0001;
  assign mem[4] = 4'b0010;
  assign mem[5] = 4'b1111;
  assign mem[6] = 4'b1011;
  assign mem[7] = 4'b1000;
  assign mem[8] = 4'b0011;
  assign mem[9] = 4'b1010;
  assign mem[10] = 4'b0110;
  assign mem[11] = 4'b1100;
  assign mem[12] = 4'b0101;
  assign mem[13] = 4'b1001;
  assign mem[14] = 4'b0000;
  assign mem[15] = 4'b0111;
  assign mem[16] = 4'b0000;
  assign mem[17] = 4'b1111;
  assign mem[18] = 4'b0111;
  assign mem[19] = 4'b0100;
  assign mem[20] = 4'b1110;
  assign mem[21] = 4'b0010;
  assign mem[22] = 4'b1101;
  assign mem[23] = 4'b0001;
  assign mem[24] = 4'b1010;
  assign mem[25] = 4'b0110;
  assign mem[26] = 4'b1100;
  assign mem[27] = 4'b1011;
  assign mem[28] = 4'b1001;
  assign mem[29] = 4'b0101;
  assign mem[30] = 4'b0011;
  assign mem[31] = 4'b1000;
  assign mem[32] = 4'b0100;
  assign mem[33] = 4'b0001;
  assign mem[34] = 4'b1110;
  assign mem[35] = 4'b1000;
  assign mem[36] = 4'b1101;
  assign mem[37] = 4'b0110;
  assign mem[38] = 4'b0010;
  assign mem[39] = 4'b1011;
  assign mem[40] = 4'b1111;
  assign mem[41] = 4'b1100;
  assign mem[42] = 4'b1001;
  assign mem[43] = 4'b0111;
  assign mem[44] = 4'b0011;
  assign mem[45] = 4'b1010;
  assign mem[46] = 4'b0101;
  assign mem[47] = 4'b0000;
  assign mem[48] = 4'b1111;
  assign mem[49] = 4'b1100;
  assign mem[50] = 4'b1000;
  assign mem[51] = 4'b0010;
  assign mem[52] = 4'b0100;
  assign mem[53] = 4'b1001;
  assign mem[54] = 4'b0001;
  assign mem[55] = 4'b0111;
  assign mem[56] = 4'b0101;
  assign mem[57] = 4'b1011;
  assign mem[58] = 4'b0011;
  assign mem[59] = 4'b1110;
  assign mem[60] = 4'b1010;
  assign mem[61] = 4'b0000;
  assign mem[62] = 4'b0110;
  assign mem[63] = 4'b1101;
  assign mem[64] = 4'b1111;
  assign mem[65] = 4'b0001;
  assign mem[66] = 4'b1000;
  assign mem[67] = 4'b1110;
  assign mem[68] = 4'b0110;
  assign mem[69] = 4'b1011;
  assign mem[70] = 4'b0011;
  assign mem[71] = 4'b0100;
  assign mem[72] = 4'b1001;
  assign mem[73] = 4'b0111;
  assign mem[74] = 4'b0010;
  assign mem[75] = 4'b1101;
  assign mem[76] = 4'b1100;
  assign mem[77] = 4'b0000;
  assign mem[78] = 4'b0101;
  assign mem[79] = 4'b1010;
  assign mem[80] = 4'b0011;
  assign mem[81] = 4'b1101;
  assign mem[82] = 4'b0100;
  assign mem[83] = 4'b0111;
  assign mem[84] = 4'b1111;
  assign mem[85] = 4'b0010;
  assign mem[86] = 4'b1000;
  assign mem[87] = 4'b1110;
  assign mem[88] = 4'b1100;
  assign mem[89] = 4'b0000;
  assign mem[90] = 4'b0001;
  assign mem[91] = 4'b1010;
  assign mem[92] = 4'b0110;
  assign mem[93] = 4'b1001;
  assign mem[94] = 4'b1011;
  assign mem[95] = 4'b0101;
  assign mem[96] = 4'b0000;
  assign mem[97] = 4'b1110;
  assign mem[98] = 4'b0111;
  assign mem[99] = 4'b1011;
  assign mem[100] = 4'b1010;
  assign mem[101] = 4'b0100;
  assign mem[102] = 4'b1101;
  assign mem[103] = 4'b0001;
  assign mem[104] = 4'b0101;
  assign mem[105] = 4'b1000;
  assign mem[106] = 4'b1100;
  assign mem[107] = 4'b0110;
  assign mem[108] = 4'b1001;
  assign mem[109] = 4'b0011;
  assign mem[110] = 4'b0010;
  assign mem[111] = 4'b1111;
  assign mem[112] = 4'b1101;
  assign mem[113] = 4'b1000;
  assign mem[114] = 4'b1010;
  assign mem[115] = 4'b0001;
  assign mem[116] = 4'b0011;
  assign mem[117] = 4'b1111;
  assign mem[118] = 4'b0100;
  assign mem[119] = 4'b0010;
  assign mem[120] = 4'b1011;
  assign mem[121] = 4'b0110;
  assign mem[122] = 4'b0111;
  assign mem[123] = 4'b1100;
  assign mem[124] = 4'b0000;
  assign mem[125] = 4'b0101;
  assign mem[126] = 4'b1110;
  assign mem[127] = 4'b1001;
  assign mem[128] = 4'b1010;
  assign mem[129] = 4'b0000;
  assign mem[130] = 4'b1001;
  assign mem[131] = 4'b1110;
  assign mem[132] = 4'b0110;
  assign mem[133] = 4'b0011;
  assign mem[134] = 4'b1111;
  assign mem[135] = 4'b0101;
  assign mem[136] = 4'b0001;
  assign mem[137] = 4'b1101;
  assign mem[138] = 4'b1100;
  assign mem[139] = 4'b0111;
  assign mem[140] = 4'b1011;
  assign mem[141] = 4'b0100;
  assign mem[142] = 4'b0010;
  assign mem[143] = 4'b1000;
  assign mem[144] = 4'b1101;
  assign mem[145] = 4'b0111;
  assign mem[146] = 4'b0000;
  assign mem[147] = 4'b1001;
  assign mem[148] = 4'b0011;
  assign mem[149] = 4'b0100;
  assign mem[150] = 4'b0110;
  assign mem[151] = 4'b1010;
  assign mem[152] = 4'b0010;
  assign mem[153] = 4'b1000;
  assign mem[154] = 4'b0101;
  assign mem[155] = 4'b1110;
  assign mem[156] = 4'b1100;
  assign mem[157] = 4'b1011;
  assign mem[158] = 4'b1111;
  assign mem[159] = 4'b0001;
  assign mem[160] = 4'b1101;
  assign mem[161] = 4'b0110;
  assign mem[162] = 4'b0100;
  assign mem[163] = 4'b1001;
  assign mem[164] = 4'b1000;
  assign mem[165] = 4'b1111;
  assign mem[166] = 4'b0011;
  assign mem[167] = 4'b0000;
  assign mem[168] = 4'b1011;
  assign mem[169] = 4'b0001;
  assign mem[170] = 4'b0010;
  assign mem[171] = 4'b1100;
  assign mem[172] = 4'b0101;
  assign mem[173] = 4'b1010;
  assign mem[174] = 4'b1110;
  assign mem[175] = 4'b0111;
  assign mem[176] = 4'b0001;
  assign mem[177] = 4'b1010;
  assign mem[178] = 4'b1101;
  assign mem[179] = 4'b0000;
  assign mem[180] = 4'b0110;
  assign mem[181] = 4'b1001;
  assign mem[182] = 4'b1000;
  assign mem[183] = 4'b0111;
  assign mem[184] = 4'b0100;
  assign mem[185] = 4'b1111;
  assign mem[186] = 4'b1110;
  assign mem[187] = 4'b0011;
  assign mem[188] = 4'b1011;
  assign mem[189] = 4'b0101;
  assign mem[190] = 4'b0010;
  assign mem[191] = 4'b1100;
  assign mem[192] = 4'b0111;
  assign mem[193] = 4'b1101;
  assign mem[194] = 4'b1110;
  assign mem[195] = 4'b0011;
  assign mem[196] = 4'b0000;
  assign mem[197] = 4'b0110;
  assign mem[198] = 4'b1001;
  assign mem[199] = 4'b1010;
  assign mem[200] = 4'b0001;
  assign mem[201] = 4'b0010;
  assign mem[202] = 4'b1000;
  assign mem[203] = 4'b0101;
  assign mem[204] = 4'b1011;
  assign mem[205] = 4'b1100;
  assign mem[206] = 4'b0100;
  assign mem[207] = 4'b1111;
  assign mem[208] = 4'b1101;
  assign mem[209] = 4'b1000;
  assign mem[210] = 4'b1011;
  assign mem[211] = 4'b0101;
  assign mem[212] = 4'b0110;
  assign mem[213] = 4'b1111;
  assign mem[214] = 4'b0000;
  assign mem[215] = 4'b0011;
  assign mem[216] = 4'b0100;
  assign mem[217] = 4'b0111;
  assign mem[218] = 4'b0010;
  assign mem[219] = 4'b1100;
  assign mem[220] = 4'b0001;
  assign mem[221] = 4'b1010;
  assign mem[222] = 4'b1110;
  assign mem[223] = 4'b1001;
  assign mem[224] = 4'b1010;
  assign mem[225] = 4'b0110;
  assign mem[226] = 4'b1001;
  assign mem[227] = 4'b0000;
  assign mem[228] = 4'b1100;
  assign mem[229] = 4'b1011;
  assign mem[230] = 4'b0111;
  assign mem[231] = 4'b1101;
  assign mem[232] = 4'b1111;
  assign mem[233] = 4'b0001;
  assign mem[234] = 4'b0011;
  assign mem[235] = 4'b1110;
  assign mem[236] = 4'b0101;
  assign mem[237] = 4'b0010;
  assign mem[238] = 4'b1000;
  assign mem[239] = 4'b0100;
  assign mem[240] = 4'b0011;
  assign mem[241] = 4'b1111;
  assign mem[242] = 4'b0000;
  assign mem[243] = 4'b0110;
  assign mem[244] = 4'b1010;
  assign mem[245] = 4'b0001;
  assign mem[246] = 4'b1101;
  assign mem[247] = 4'b1000;
  assign mem[248] = 4'b1001;
  assign mem[249] = 4'b0100;
  assign mem[250] = 4'b0101;
  assign mem[251] = 4'b1011;
  assign mem[252] = 4'b1100;
  assign mem[253] = 4'b0111;
  assign mem[254] = 4'b0010;
  assign mem[255] = 4'b1110;
  assign mem[256] = 4'b0010;
  assign mem[257] = 4'b1100;
  assign mem[258] = 4'b0100;
  assign mem[259] = 4'b0001;
  assign mem[260] = 4'b0111;
  assign mem[261] = 4'b1010;
  assign mem[262] = 4'b1011;
  assign mem[263] = 4'b0110;
  assign mem[264] = 4'b1000;
  assign mem[265] = 4'b0101;
  assign mem[266] = 4'b0011;
  assign mem[267] = 4'b1111;
  assign mem[268] = 4'b1101;
  assign mem[269] = 4'b0000;
  assign mem[270] = 4'b1110;
  assign mem[271] = 4'b1001;
  assign mem[272] = 4'b1110;
  assign mem[273] = 4'b1011;
  assign mem[274] = 4'b0010;
  assign mem[275] = 4'b1100;
  assign mem[276] = 4'b0100;
  assign mem[277] = 4'b0111;
  assign mem[278] = 4'b1101;
  assign mem[279] = 4'b0001;
  assign mem[280] = 4'b0101;
  assign mem[281] = 4'b0000;
  assign mem[282] = 4'b1111;
  assign mem[283] = 4'b1010;
  assign mem[284] = 4'b0011;
  assign mem[285] = 4'b1001;
  assign mem[286] = 4'b1000;
  assign mem[287] = 4'b0110;
  assign mem[288] = 4'b0100;
  assign mem[289] = 4'b0010;
  assign mem[290] = 4'b0001;
  assign mem[291] = 4'b1011;
  assign mem[292] = 4'b1010;
  assign mem[293] = 4'b1101;
  assign mem[294] = 4'b0111;
  assign mem[295] = 4'b1000;
  assign mem[296] = 4'b1111;
  assign mem[297] = 4'b1001;
  assign mem[298] = 4'b1100;
  assign mem[299] = 4'b0101;
  assign mem[300] = 4'b0110;
  assign mem[301] = 4'b0011;
  assign mem[302] = 4'b0000;
  assign mem[303] = 4'b1110;
  assign mem[304] = 4'b1011;
  assign mem[305] = 4'b1000;
  assign mem[306] = 4'b1100;
  assign mem[307] = 4'b0111;
  assign mem[308] = 4'b0001;
  assign mem[309] = 4'b1110;
  assign mem[310] = 4'b0010;
  assign mem[311] = 4'b1101;
  assign mem[312] = 4'b0110;
  assign mem[313] = 4'b1111;
  assign mem[314] = 4'b0000;
  assign mem[315] = 4'b1001;
  assign mem[316] = 4'b1010;
  assign mem[317] = 4'b0100;
  assign mem[318] = 4'b0101;
  assign mem[319] = 4'b0011;
  assign mem[320] = 4'b1100;
  assign mem[321] = 4'b0001;
  assign mem[322] = 4'b1010;
  assign mem[323] = 4'b1111;
  assign mem[324] = 4'b1001;
  assign mem[325] = 4'b0010;
  assign mem[326] = 4'b0110;
  assign mem[327] = 4'b1000;
  assign mem[328] = 4'b0000;
  assign mem[329] = 4'b1101;
  assign mem[330] = 4'b0011;
  assign mem[331] = 4'b0100;
  assign mem[332] = 4'b1110;
  assign mem[333] = 4'b0111;
  assign mem[334] = 4'b0101;
  assign mem[335] = 4'b1011;
  assign mem[336] = 4'b1010;
  assign mem[337] = 4'b1111;
  assign mem[338] = 4'b0100;
  assign mem[339] = 4'b0010;
  assign mem[340] = 4'b0111;
  assign mem[341] = 4'b1100;
  assign mem[342] = 4'b1001;
  assign mem[343] = 4'b0101;
  assign mem[344] = 4'b0110;
  assign mem[345] = 4'b0001;
  assign mem[346] = 4'b1101;
  assign mem[347] = 4'b1110;
  assign mem[348] = 4'b0000;
  assign mem[349] = 4'b1011;
  assign mem[350] = 4'b0011;
  assign mem[351] = 4'b1000;
  assign mem[352] = 4'b1001;
  assign mem[353] = 4'b1110;
  assign mem[354] = 4'b1111;
  assign mem[355] = 4'b0101;
  assign mem[356] = 4'b0010;
  assign mem[357] = 4'b1000;
  assign mem[358] = 4'b1100;
  assign mem[359] = 4'b0011;
  assign mem[360] = 4'b0111;
  assign mem[361] = 4'b0000;
  assign mem[362] = 4'b0100;
  assign mem[363] = 4'b1010;
  assign mem[364] = 4'b0001;
  assign mem[365] = 4'b1101;
  assign mem[366] = 4'b1011;
  assign mem[367] = 4'b0110;
  assign mem[368] = 4'b0100;
  assign mem[369] = 4'b0011;
  assign mem[370] = 4'b0010;
  assign mem[371] = 4'b1100;
  assign mem[372] = 4'b1001;
  assign mem[373] = 4'b0101;
  assign mem[374] = 4'b1111;
  assign mem[375] = 4'b1010;
  assign mem[376] = 4'b1011;
  assign mem[377] = 4'b1110;
  assign mem[378] = 4'b0001;
  assign mem[379] = 4'b0111;
  assign mem[380] = 4'b0110;
  assign mem[381] = 4'b0000;
  assign mem[382] = 4'b1000;
  assign mem[383] = 4'b1101;
  assign mem[384] = 4'b0100;
  assign mem[385] = 4'b1011;
  assign mem[386] = 4'b0010;
  assign mem[387] = 4'b1110;
  assign mem[388] = 4'b1111;
  assign mem[389] = 4'b0000;
  assign mem[390] = 4'b1000;
  assign mem[391] = 4'b1101;
  assign mem[392] = 4'b0011;
  assign mem[393] = 4'b1100;
  assign mem[394] = 4'b1001;
  assign mem[395] = 4'b0111;
  assign mem[396] = 4'b0101;
  assign mem[397] = 4'b1010;
  assign mem[398] = 4'b0110;
  assign mem[399] = 4'b0001;
  assign mem[400] = 4'b1101;
  assign mem[401] = 4'b0000;
  assign mem[402] = 4'b1011;
  assign mem[403] = 4'b0111;
  assign mem[404] = 4'b0100;
  assign mem[405] = 4'b1001;
  assign mem[406] = 4'b0001;
  assign mem[407] = 4'b1010;
  assign mem[408] = 4'b1110;
  assign mem[409] = 4'b0011;
  assign mem[410] = 4'b0101;
  assign mem[411] = 4'b1100;
  assign mem[412] = 4'b0010;
  assign mem[413] = 4'b1111;
  assign mem[414] = 4'b1000;
  assign mem[415] = 4'b0110;
  assign mem[416] = 4'b0001;
  assign mem[417] = 4'b0100;
  assign mem[418] = 4'b1011;
  assign mem[419] = 4'b1101;
  assign mem[420] = 4'b1100;
  assign mem[421] = 4'b0011;
  assign mem[422] = 4'b0111;
  assign mem[423] = 4'b1110;
  assign mem[424] = 4'b1010;
  assign mem[425] = 4'b1111;
  assign mem[426] = 4'b0110;
  assign mem[427] = 4'b1000;
  assign mem[428] = 4'b0000;
  assign mem[429] = 4'b0101;
  assign mem[430] = 4'b1001;
  assign mem[431] = 4'b0010;
  assign mem[432] = 4'b0110;
  assign mem[433] = 4'b1011;
  assign mem[434] = 4'b1101;
  assign mem[435] = 4'b1000;
  assign mem[436] = 4'b0001;
  assign mem[437] = 4'b0100;
  assign mem[438] = 4'b1010;
  assign mem[439] = 4'b0111;
  assign mem[440] = 4'b1001;
  assign mem[441] = 4'b0101;
  assign mem[442] = 4'b0000;
  assign mem[443] = 4'b1111;
  assign mem[444] = 4'b1110;
  assign mem[445] = 4'b0010;
  assign mem[446] = 4'b0011;
  assign mem[447] = 4'b1100;
  assign mem[448] = 4'b1101;
  assign mem[449] = 4'b0010;
  assign mem[450] = 4'b1000;
  assign mem[451] = 4'b0100;
  assign mem[452] = 4'b0110;
  assign mem[453] = 4'b1111;
  assign mem[454] = 4'b1011;
  assign mem[455] = 4'b0001;
  assign mem[456] = 4'b1010;
  assign mem[457] = 4'b1001;
  assign mem[458] = 4'b0011;
  assign mem[459] = 4'b1110;
  assign mem[460] = 4'b0101;
  assign mem[461] = 4'b0000;
  assign mem[462] = 4'b1100;
  assign mem[463] = 4'b0111;
  assign mem[464] = 4'b0001;
  assign mem[465] = 4'b1111;
  assign mem[466] = 4'b1101;
  assign mem[467] = 4'b1000;
  assign mem[468] = 4'b1010;
  assign mem[469] = 4'b0011;
  assign mem[470] = 4'b0111;
  assign mem[471] = 4'b0100;
  assign mem[472] = 4'b1100;
  assign mem[473] = 4'b0101;
  assign mem[474] = 4'b0110;
  assign mem[475] = 4'b1011;
  assign mem[476] = 4'b0000;
  assign mem[477] = 4'b1110;
  assign mem[478] = 4'b1001;
  assign mem[479] = 4'b0010;
  assign mem[480] = 4'b0111;
  assign mem[481] = 4'b1011;
  assign mem[482] = 4'b0100;
  assign mem[483] = 4'b0001;
  assign mem[484] = 4'b1001;
  assign mem[485] = 4'b1100;
  assign mem[486] = 4'b1110;
  assign mem[487] = 4'b0010;
  assign mem[488] = 4'b0000;
  assign mem[489] = 4'b0110;
  assign mem[490] = 4'b1010;
  assign mem[491] = 4'b1101;
  assign mem[492] = 4'b1111;
  assign mem[493] = 4'b0011;
  assign mem[494] = 4'b0101;
  assign mem[495] = 4'b1000;
  assign mem[496] = 4'b0010;
  assign mem[497] = 4'b0001;
  assign mem[498] = 4'b1110;
  assign mem[499] = 4'b0111;
  assign mem[500] = 4'b0100;
  assign mem[501] = 4'b1010;
  assign mem[502] = 4'b1000;
  assign mem[503] = 4'b1101;
  assign mem[504] = 4'b1111;
  assign mem[505] = 4'b1100;
  assign mem[506] = 4'b1001;
  assign mem[507] = 4'b0000;
  assign mem[508] = 4'b0011;
  assign mem[509] = 4'b0101;
  assign mem[510] = 4'b0110;
  assign mem[511] = 4'b1011;


  // Combinational ROM read block
  always@(*)
  begin
    data_out_t <= mem[addr];
  end

  // Output register assignment
  assign data_out = data_out_t;

endmodule



//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Sun Mar 21 12:44:04 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    des_check_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module des_check_core_core_fsm (
  clk, rst, fsm_output
);
  input clk;
  input rst;
  output [16:0] fsm_output;
  reg [16:0] fsm_output;


  // FSM State Type Declaration for des_check_core_core_fsm_1
  parameter
    main_C_0 = 5'd0,
    main_C_1 = 5'd1,
    main_C_2 = 5'd2,
    main_C_3 = 5'd3,
    main_C_4 = 5'd4,
    main_C_5 = 5'd5,
    main_C_6 = 5'd6,
    main_C_7 = 5'd7,
    main_C_8 = 5'd8,
    main_C_9 = 5'd9,
    main_C_10 = 5'd10,
    main_C_11 = 5'd11,
    main_C_12 = 5'd12,
    main_C_13 = 5'd13,
    main_C_14 = 5'd14,
    main_C_15 = 5'd15,
    main_C_16 = 5'd16;

  reg [4:0] state_var;
  reg [4:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : des_check_core_core_fsm_1
    case (state_var)
      main_C_1 : begin
        fsm_output = 17'b00000000000000010;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 17'b00000000000000100;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 17'b00000000000001000;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 17'b00000000000010000;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 17'b00000000000100000;
        state_var_NS = main_C_6;
      end
      main_C_6 : begin
        fsm_output = 17'b00000000001000000;
        state_var_NS = main_C_7;
      end
      main_C_7 : begin
        fsm_output = 17'b00000000010000000;
        state_var_NS = main_C_8;
      end
      main_C_8 : begin
        fsm_output = 17'b00000000100000000;
        state_var_NS = main_C_9;
      end
      main_C_9 : begin
        fsm_output = 17'b00000001000000000;
        state_var_NS = main_C_10;
      end
      main_C_10 : begin
        fsm_output = 17'b00000010000000000;
        state_var_NS = main_C_11;
      end
      main_C_11 : begin
        fsm_output = 17'b00000100000000000;
        state_var_NS = main_C_12;
      end
      main_C_12 : begin
        fsm_output = 17'b00001000000000000;
        state_var_NS = main_C_13;
      end
      main_C_13 : begin
        fsm_output = 17'b00010000000000000;
        state_var_NS = main_C_14;
      end
      main_C_14 : begin
        fsm_output = 17'b00100000000000000;
        state_var_NS = main_C_15;
      end
      main_C_15 : begin
        fsm_output = 17'b01000000000000000;
        state_var_NS = main_C_16;
      end
      main_C_16 : begin
        fsm_output = 17'b10000000000000000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 17'b00000000000000001;
        state_var_NS = main_C_1;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    des_check_core
// ------------------------------------------------------------------


module des_check_core (
  clk, rst, input_rsc_dat, input_rsc_triosy_lz, key_rsc_dat, key_rsc_triosy_lz, return_rsc_dat,
      return_rsc_triosy_lz
);
  input clk;
  input rst;
  input [63:0] input_rsc_dat;
  output input_rsc_triosy_lz;
  input [63:0] key_rsc_dat;
  output key_rsc_triosy_lz;
  output [63:0] return_rsc_dat;
  output return_rsc_triosy_lz;


  // Interconnect Declarations
  wire [63:0] input_rsci_idat;
  wire [63:0] key_rsci_idat;
  reg return_rsc_triosy_obj_ld;
  reg return_rsci_idat_63;
  reg return_rsci_idat_62;
  reg return_rsci_idat_61;
  reg return_rsci_idat_60;
  reg return_rsci_idat_59;
  reg return_rsci_idat_58;
  reg return_rsci_idat_57;
  reg return_rsci_idat_56;
  reg return_rsci_idat_55;
  reg return_rsci_idat_54;
  reg return_rsci_idat_53;
  reg return_rsci_idat_52;
  reg return_rsci_idat_51;
  reg return_rsci_idat_50;
  reg return_rsci_idat_49;
  reg return_rsci_idat_48;
  reg return_rsci_idat_47;
  reg return_rsci_idat_46;
  reg return_rsci_idat_45;
  reg return_rsci_idat_44;
  reg return_rsci_idat_43;
  reg return_rsci_idat_42;
  reg return_rsci_idat_41;
  reg return_rsci_idat_40;
  reg return_rsci_idat_39;
  reg return_rsci_idat_38;
  reg return_rsci_idat_37;
  reg return_rsci_idat_36;
  reg return_rsci_idat_35;
  reg return_rsci_idat_34;
  reg return_rsci_idat_33;
  reg return_rsci_idat_32;
  reg return_rsci_idat_31;
  reg return_rsci_idat_30;
  reg return_rsci_idat_29;
  reg return_rsci_idat_28;
  reg return_rsci_idat_27;
  reg return_rsci_idat_26;
  reg return_rsci_idat_25;
  reg return_rsci_idat_24;
  reg return_rsci_idat_23;
  reg return_rsci_idat_22;
  reg return_rsci_idat_21;
  reg return_rsci_idat_20;
  reg return_rsci_idat_19;
  reg return_rsci_idat_18;
  reg return_rsci_idat_17;
  reg return_rsci_idat_16;
  reg return_rsci_idat_15;
  reg return_rsci_idat_14;
  reg return_rsci_idat_13;
  reg return_rsci_idat_12;
  reg return_rsci_idat_11;
  reg return_rsci_idat_10;
  reg return_rsci_idat_9;
  reg return_rsci_idat_8;
  reg return_rsci_idat_7;
  reg return_rsci_idat_6;
  reg return_rsci_idat_5;
  reg return_rsci_idat_4;
  reg return_rsci_idat_3;
  reg return_rsci_idat_2;
  reg return_rsci_idat_1;
  reg return_rsci_idat_0;
  wire [16:0] fsm_output;
  reg reg_input_rsc_triosy_obj_ld_cse;
  wire [3:0] operator_8_false_1_read_rom_S_rom_map_1_6_itm;
  wire [3:0] operator_8_false_1_read_rom_S_rom_map_1_5_itm;
  wire [3:0] operator_8_false_1_read_rom_S_rom_map_1_2_itm;
  wire [3:0] operator_8_false_1_read_rom_S_rom_map_1_itm;
  wire [3:0] operator_8_false_1_read_rom_S_rom_map_1_1_itm;
  wire [3:0] operator_8_false_1_read_rom_S_rom_map_1_4_itm;
  wire [3:0] operator_8_false_1_read_rom_S_rom_map_1_3_itm;
  wire [3:0] operator_8_false_1_read_rom_S_rom_map_1_7_itm;
  wire [3:0] operator_8_false_1_read_rom_S_rom_map_1_14_itm;
  wire [3:0] operator_8_false_1_read_rom_S_rom_map_1_13_itm;
  wire [3:0] operator_8_false_1_read_rom_S_rom_map_1_10_itm;
  wire [3:0] operator_8_false_1_read_rom_S_rom_map_1_8_itm;
  wire [3:0] operator_8_false_1_read_rom_S_rom_map_1_9_itm;
  wire [3:0] operator_8_false_1_read_rom_S_rom_map_1_12_itm;
  wire [3:0] operator_8_false_1_read_rom_S_rom_map_1_11_itm;
  wire [3:0] operator_8_false_1_read_rom_S_rom_map_1_15_itm;
  reg [63:0] input_sva;
  reg [62:0] key_io_read_key_rsc_cse_63_1_sva;
  reg [3:0] s_output_1_19_16_19_sva;
  reg [3:0] s_output_1_3_0_23_sva;
  reg [3:0] s_output_1_19_16_34_sva;
  reg [3:0] s_output_1_3_0_38_sva;
  reg [3:0] s_output_1_19_16_49_sva;
  reg [3:0] s_output_1_3_0_53_sva;
  reg [3:0] s_output_1_19_16_4_sva;
  reg [3:0] s_output_1_3_0_8_sva;
  reg R_15_1_sva;
  reg R_16_1_sva;
  reg R_14_1_sva;
  reg R_17_1_sva;
  reg R_13_1_sva;
  reg R_18_1_sva;
  reg R_12_1_sva;
  reg R_19_1_sva;
  reg R_11_1_sva;
  reg R_20_1_sva;
  reg R_10_1_sva;
  reg R_21_1_sva;
  reg R_9_1_sva;
  reg R_22_1_sva;
  reg R_8_1_sva;
  reg R_23_1_sva;
  reg R_7_1_sva;
  reg R_24_1_sva;
  reg R_6_1_sva;
  reg R_25_1_sva;
  reg R_5_1_sva;
  reg R_26_1_sva;
  reg R_4_1_sva;
  reg R_27_1_sva;
  reg R_3_1_sva;
  reg R_28_1_sva;
  reg R_2_1_sva;
  reg R_29_1_sva;
  reg R_1_1_sva;
  reg R_30_1_sva;
  reg R_0_1_sva;
  reg R_31_1_sva;
  reg [3:0] s_output_1_19_16_20_sva;
  reg [3:0] s_output_1_3_0_24_sva;
  reg [3:0] s_output_1_19_16_35_sva;
  reg [3:0] s_output_1_3_0_39_sva;
  reg [3:0] s_output_1_19_16_50_sva;
  reg [3:0] s_output_1_3_0_54_sva;
  reg [3:0] s_output_1_19_16_5_sva;
  reg [3:0] s_output_1_3_0_9_sva;
  reg R_15_3_sva;
  reg R_16_3_sva;
  reg R_14_3_sva;
  reg R_17_3_sva;
  reg R_13_3_sva;
  reg R_18_3_sva;
  reg R_12_3_sva;
  reg R_19_3_sva;
  reg R_11_3_sva;
  reg R_20_3_sva;
  reg R_10_3_sva;
  reg R_21_3_sva;
  reg R_9_3_sva;
  reg R_22_3_sva;
  reg R_8_3_sva;
  reg R_23_3_sva;
  reg R_7_3_sva;
  reg R_24_3_sva;
  reg R_6_3_sva;
  reg R_25_3_sva;
  reg R_5_3_sva;
  reg R_26_3_sva;
  reg R_4_3_sva;
  reg R_27_3_sva;
  reg R_3_3_sva;
  reg R_28_3_sva;
  reg R_2_3_sva;
  reg R_29_3_sva;
  reg R_1_3_sva;
  reg R_30_3_sva;
  reg R_0_3_sva;
  reg R_31_3_sva;
  reg R_15_4_sva;
  reg R_16_4_sva;
  reg R_14_4_sva;
  reg R_17_4_sva;
  reg R_13_4_sva;
  reg R_18_4_sva;
  reg R_12_4_sva;
  reg R_19_4_sva;
  reg R_11_4_sva;
  reg R_20_4_sva;
  reg R_10_4_sva;
  reg R_21_4_sva;
  reg R_9_4_sva;
  reg R_22_4_sva;
  reg R_8_4_sva;
  reg R_23_4_sva;
  reg R_7_4_sva;
  reg R_24_4_sva;
  reg R_6_4_sva;
  reg R_25_4_sva;
  reg R_5_4_sva;
  reg R_26_4_sva;
  reg R_4_4_sva;
  reg R_27_4_sva;
  reg R_3_4_sva;
  reg R_28_4_sva;
  reg R_2_4_sva;
  reg R_29_4_sva;
  reg R_1_4_sva;
  reg R_30_4_sva;
  reg R_0_4_sva;
  reg R_31_4_sva;
  reg R_15_5_sva;
  reg R_16_5_sva;
  reg R_14_5_sva;
  reg R_17_5_sva;
  reg R_13_5_sva;
  reg R_18_5_sva;
  reg R_12_5_sva;
  reg R_19_5_sva;
  reg R_11_5_sva;
  reg R_20_5_sva;
  reg R_10_5_sva;
  reg R_21_5_sva;
  reg R_9_5_sva;
  reg R_22_5_sva;
  reg R_8_5_sva;
  reg R_23_5_sva;
  reg R_7_5_sva;
  reg R_24_5_sva;
  reg R_6_5_sva;
  reg R_25_5_sva;
  reg R_5_5_sva;
  reg R_26_5_sva;
  reg R_4_5_sva;
  reg R_27_5_sva;
  reg R_3_5_sva;
  reg R_28_5_sva;
  reg R_2_5_sva;
  reg R_29_5_sva;
  reg R_1_5_sva;
  reg R_30_5_sva;
  reg R_0_5_sva;
  reg R_31_5_sva;
  reg R_15_6_sva;
  reg R_16_6_sva;
  reg R_14_6_sva;
  reg R_17_6_sva;
  reg R_13_6_sva;
  reg R_18_6_sva;
  reg R_12_6_sva;
  reg R_19_6_sva;
  reg R_11_6_sva;
  reg R_20_6_sva;
  reg R_10_6_sva;
  reg R_21_6_sva;
  reg R_9_6_sva;
  reg R_22_6_sva;
  reg R_8_6_sva;
  reg R_23_6_sva;
  reg R_7_6_sva;
  reg R_24_6_sva;
  reg R_6_6_sva;
  reg R_25_6_sva;
  reg R_5_6_sva;
  reg R_26_6_sva;
  reg R_4_6_sva;
  reg R_27_6_sva;
  reg R_3_6_sva;
  reg R_28_6_sva;
  reg R_2_6_sva;
  reg R_29_6_sva;
  reg R_1_6_sva;
  reg R_30_6_sva;
  reg R_0_6_sva;
  reg R_31_6_sva;
  reg R_15_7_sva;
  reg R_16_7_sva;
  reg R_14_7_sva;
  reg R_17_7_sva;
  reg R_13_7_sva;
  reg R_18_7_sva;
  reg R_12_7_sva;
  reg R_19_7_sva;
  reg R_11_7_sva;
  reg R_20_7_sva;
  reg R_10_7_sva;
  reg R_21_7_sva;
  reg R_9_7_sva;
  reg R_22_7_sva;
  reg R_8_7_sva;
  reg R_23_7_sva;
  reg R_7_7_sva;
  reg R_24_7_sva;
  reg R_6_7_sva;
  reg R_25_7_sva;
  reg R_5_7_sva;
  reg R_26_7_sva;
  reg R_4_7_sva;
  reg R_27_7_sva;
  reg R_3_7_sva;
  reg R_28_7_sva;
  reg R_2_7_sva;
  reg R_29_7_sva;
  reg R_1_7_sva;
  reg R_30_7_sva;
  reg R_0_7_sva;
  reg R_31_7_sva;
  reg R_15_8_sva;
  reg R_16_8_sva;
  reg R_14_8_sva;
  reg R_17_8_sva;
  reg R_13_8_sva;
  reg R_18_8_sva;
  reg R_12_8_sva;
  reg R_19_8_sva;
  reg R_11_8_sva;
  reg R_20_8_sva;
  reg R_10_8_sva;
  reg R_21_8_sva;
  reg R_9_8_sva;
  reg R_22_8_sva;
  reg R_8_8_sva;
  reg R_23_8_sva;
  reg R_7_8_sva;
  reg R_24_8_sva;
  reg R_6_8_sva;
  reg R_25_8_sva;
  reg R_5_8_sva;
  reg R_26_8_sva;
  reg R_4_8_sva;
  reg R_27_8_sva;
  reg R_3_8_sva;
  reg R_28_8_sva;
  reg R_2_8_sva;
  reg R_29_8_sva;
  reg R_1_8_sva;
  reg R_30_8_sva;
  reg R_0_8_sva;
  reg R_31_8_sva;
  reg R_15_9_sva;
  reg R_16_9_sva;
  reg R_14_9_sva;
  reg R_17_9_sva;
  reg R_13_9_sva;
  reg R_18_9_sva;
  reg R_12_9_sva;
  reg R_19_9_sva;
  reg R_11_9_sva;
  reg R_20_9_sva;
  reg R_10_9_sva;
  reg R_21_9_sva;
  reg R_9_9_sva;
  reg R_22_9_sva;
  reg R_8_9_sva;
  reg R_23_9_sva;
  reg R_7_9_sva;
  reg R_24_9_sva;
  reg R_6_9_sva;
  reg R_25_9_sva;
  reg R_5_9_sva;
  reg R_26_9_sva;
  reg R_4_9_sva;
  reg R_27_9_sva;
  reg R_3_9_sva;
  reg R_28_9_sva;
  reg R_2_9_sva;
  reg R_29_9_sva;
  reg R_1_9_sva;
  reg R_30_9_sva;
  reg R_0_9_sva;
  reg R_31_9_sva;
  reg R_15_10_sva;
  reg R_16_10_sva;
  reg R_14_10_sva;
  reg R_17_10_sva;
  reg R_13_10_sva;
  reg R_18_10_sva;
  reg R_12_10_sva;
  reg R_19_10_sva;
  reg R_11_10_sva;
  reg R_20_10_sva;
  reg R_10_10_sva;
  reg R_21_10_sva;
  reg R_9_10_sva;
  reg R_22_10_sva;
  reg R_8_10_sva;
  reg R_23_10_sva;
  reg R_7_10_sva;
  reg R_24_10_sva;
  reg R_6_10_sva;
  reg R_25_10_sva;
  reg R_5_10_sva;
  reg R_26_10_sva;
  reg R_4_10_sva;
  reg R_27_10_sva;
  reg R_3_10_sva;
  reg R_28_10_sva;
  reg R_2_10_sva;
  reg R_29_10_sva;
  reg R_1_10_sva;
  reg R_30_10_sva;
  reg R_0_10_sva;
  reg R_31_10_sva;
  reg R_15_11_sva;
  reg R_16_11_sva;
  reg R_14_11_sva;
  reg R_17_11_sva;
  reg R_13_11_sva;
  reg R_18_11_sva;
  reg R_12_11_sva;
  reg R_19_11_sva;
  reg R_11_11_sva;
  reg R_20_11_sva;
  reg R_10_11_sva;
  reg R_21_11_sva;
  reg R_9_11_sva;
  reg R_22_11_sva;
  reg R_8_11_sva;
  reg R_23_11_sva;
  reg R_7_11_sva;
  reg R_24_11_sva;
  reg R_6_11_sva;
  reg R_25_11_sva;
  reg R_5_11_sva;
  reg R_26_11_sva;
  reg R_4_11_sva;
  reg R_27_11_sva;
  reg R_3_11_sva;
  reg R_28_11_sva;
  reg R_2_11_sva;
  reg R_29_11_sva;
  reg R_1_11_sva;
  reg R_30_11_sva;
  reg R_0_11_sva;
  reg R_31_11_sva;
  reg R_15_12_sva;
  reg R_16_12_sva;
  reg R_14_12_sva;
  reg R_17_12_sva;
  reg R_13_12_sva;
  reg R_18_12_sva;
  reg R_12_12_sva;
  reg R_19_12_sva;
  reg R_11_12_sva;
  reg R_20_12_sva;
  reg R_10_12_sva;
  reg R_21_12_sva;
  reg R_9_12_sva;
  reg R_22_12_sva;
  reg R_8_12_sva;
  reg R_23_12_sva;
  reg R_7_12_sva;
  reg R_24_12_sva;
  reg R_6_12_sva;
  reg R_25_12_sva;
  reg R_5_12_sva;
  reg R_26_12_sva;
  reg R_4_12_sva;
  reg R_27_12_sva;
  reg R_3_12_sva;
  reg R_28_12_sva;
  reg R_2_12_sva;
  reg R_29_12_sva;
  reg R_1_12_sva;
  reg R_30_12_sva;
  reg R_0_12_sva;
  reg R_31_12_sva;
  reg R_15_13_sva;
  reg R_16_13_sva;
  reg R_14_13_sva;
  reg R_17_13_sva;
  reg R_13_13_sva;
  reg R_18_13_sva;
  reg R_12_13_sva;
  reg R_19_13_sva;
  reg R_11_13_sva;
  reg R_20_13_sva;
  reg R_10_13_sva;
  reg R_21_13_sva;
  reg R_9_13_sva;
  reg R_22_13_sva;
  reg R_8_13_sva;
  reg R_23_13_sva;
  reg R_7_13_sva;
  reg R_24_13_sva;
  reg R_6_13_sva;
  reg R_25_13_sva;
  reg R_5_13_sva;
  reg R_26_13_sva;
  reg R_4_13_sva;
  reg R_27_13_sva;
  reg R_3_13_sva;
  reg R_28_13_sva;
  reg R_2_13_sva;
  reg R_29_13_sva;
  reg R_1_13_sva;
  reg R_30_13_sva;
  reg R_0_13_sva;
  reg R_31_13_sva;
  reg R_15_14_sva;
  reg R_16_14_sva;
  reg R_14_14_sva;
  reg R_17_14_sva;
  reg R_13_14_sva;
  reg R_18_14_sva;
  reg R_12_14_sva;
  reg R_19_14_sva;
  reg R_11_14_sva;
  reg R_20_14_sva;
  reg R_10_14_sva;
  reg R_21_14_sva;
  reg R_9_14_sva;
  reg R_22_14_sva;
  reg R_8_14_sva;
  reg R_23_14_sva;
  reg R_7_14_sva;
  reg R_24_14_sva;
  reg R_6_14_sva;
  reg R_25_14_sva;
  reg R_5_14_sva;
  reg R_26_14_sva;
  reg R_4_14_sva;
  reg R_27_14_sva;
  reg R_3_14_sva;
  reg R_28_14_sva;
  reg R_2_14_sva;
  reg R_29_14_sva;
  reg R_1_14_sva;
  reg R_30_14_sva;
  reg R_0_14_sva;
  reg R_31_14_sva;
  reg R_15_15_sva;
  reg R_16_15_sva;
  reg R_14_15_sva;
  reg R_17_15_sva;
  reg R_13_15_sva;
  reg R_18_15_sva;
  reg R_12_15_sva;
  reg R_19_15_sva;
  reg R_11_15_sva;
  reg R_20_15_sva;
  reg R_10_15_sva;
  reg R_21_15_sva;
  reg R_9_15_sva;
  reg R_22_15_sva;
  reg R_8_15_sva;
  reg R_23_15_sva;
  reg R_7_15_sva;
  reg R_24_15_sva;
  reg R_6_15_sva;
  reg R_25_15_sva;
  reg R_5_15_sva;
  reg R_26_15_sva;
  reg R_4_15_sva;
  reg R_27_15_sva;
  reg R_3_15_sva;
  reg R_28_15_sva;
  reg R_2_15_sva;
  reg R_29_15_sva;
  reg R_1_15_sva;
  reg R_30_15_sva;
  reg R_0_15_sva;
  reg R_31_15_sva;
  wire [3:0] s_output_1_19_16_6_sva_1;
  wire [3:0] s_output_1_3_0_55_sva_1;
  wire [3:0] s_output_1_19_16_36_sva_1;
  wire [3:0] s_output_1_19_16_21_sva_1;
  wire [3:0] s_output_1_3_0_25_sva_1;
  wire [3:0] s_output_1_19_16_51_sva_1;
  wire [3:0] s_output_1_3_0_40_sva_1;
  wire [3:0] s_output_1_3_0_10_sva_1;
  wire [3:0] s_output_1_19_16_7_sva_1;
  wire [3:0] s_output_1_3_0_56_sva_1;
  wire [3:0] s_output_1_19_16_37_sva_1;
  wire [3:0] s_output_1_19_16_22_sva_1;
  wire [3:0] s_output_1_3_0_26_sva_1;
  wire [3:0] s_output_1_19_16_52_sva_1;
  wire [3:0] s_output_1_3_0_41_sva_1;
  wire [3:0] s_output_1_3_0_11_sva_1;
  wire [3:0] s_output_1_19_16_8_sva_1;
  wire [3:0] s_output_1_3_0_57_sva_1;
  wire [3:0] s_output_1_19_16_38_sva_1;
  wire [3:0] s_output_1_19_16_23_sva_1;
  wire [3:0] s_output_1_3_0_27_sva_1;
  wire [3:0] s_output_1_19_16_53_sva_1;
  wire [3:0] s_output_1_3_0_42_sva_1;
  wire [3:0] s_output_1_3_0_12_sva_1;
  wire [3:0] s_output_1_19_16_9_sva_1;
  wire [3:0] s_output_1_3_0_58_sva_1;
  wire [3:0] s_output_1_19_16_39_sva_1;
  wire [3:0] s_output_1_19_16_24_sva_1;
  wire [3:0] s_output_1_3_0_28_sva_1;
  wire [3:0] s_output_1_19_16_54_sva_1;
  wire [3:0] s_output_1_3_0_43_sva_1;
  wire [3:0] s_output_1_3_0_13_sva_1;
  wire [3:0] s_output_1_19_16_10_sva_1;
  wire [3:0] s_output_1_3_0_59_sva_1;
  wire [3:0] s_output_1_19_16_40_sva_1;
  wire [3:0] s_output_1_19_16_25_sva_1;
  wire [3:0] s_output_1_3_0_29_sva_1;
  wire [3:0] s_output_1_19_16_55_sva_1;
  wire [3:0] s_output_1_3_0_44_sva_1;
  wire [3:0] s_output_1_3_0_14_sva_1;
  wire [3:0] s_output_1_19_16_11_sva_1;
  wire [3:0] s_output_1_3_0_60_sva_1;
  wire [3:0] s_output_1_19_16_41_sva_1;
  wire [3:0] s_output_1_19_16_26_sva_1;
  wire [3:0] s_output_1_3_0_30_sva_1;
  wire [3:0] s_output_1_19_16_56_sva_1;
  wire [3:0] s_output_1_3_0_45_sva_1;
  wire [3:0] s_output_1_3_0_15_sva_1;
  wire [3:0] s_output_1_19_16_12_sva_1;
  wire [3:0] s_output_1_3_0_61_sva_1;
  wire [3:0] s_output_1_19_16_42_sva_1;
  wire [3:0] s_output_1_19_16_27_sva_1;
  wire [3:0] s_output_1_3_0_31_sva_1;
  wire [3:0] s_output_1_19_16_57_sva_1;
  wire [3:0] s_output_1_3_0_46_sva_1;
  wire [3:0] s_output_1_3_0_16_sva_1;
  wire [3:0] s_output_1_19_16_13_sva_1;
  wire [3:0] s_output_1_3_0_62_sva_1;
  wire [3:0] s_output_1_19_16_43_sva_1;
  wire [3:0] s_output_1_19_16_28_sva_1;
  wire [3:0] s_output_1_3_0_32_sva_1;
  wire [3:0] s_output_1_19_16_58_sva_1;
  wire [3:0] s_output_1_3_0_47_sva_1;
  wire [3:0] s_output_1_3_0_17_sva_1;
  wire [3:0] s_output_1_19_16_14_sva_1;
  wire [3:0] s_output_1_3_0_63_sva_1;
  wire [3:0] s_output_1_19_16_44_sva_1;
  wire [3:0] s_output_1_19_16_29_sva_1;
  wire [3:0] s_output_1_3_0_33_sva_1;
  wire [3:0] s_output_1_19_16_59_sva_1;
  wire [3:0] s_output_1_3_0_48_sva_1;
  wire [3:0] s_output_1_3_0_18_sva_1;
  wire [3:0] s_output_1_19_16_15_sva_1;
  wire [3:0] s_output_1_3_0_64_sva_1;
  wire [3:0] s_output_1_19_16_45_sva_1;
  wire [3:0] s_output_1_19_16_30_sva_1;
  wire [3:0] s_output_1_3_0_34_sva_1;
  wire [3:0] s_output_1_19_16_60_sva_1;
  wire [3:0] s_output_1_3_0_49_sva_1;
  wire [3:0] s_output_1_3_0_19_sva_1;
  wire [3:0] s_output_1_19_16_16_sva_1;
  wire [3:0] s_output_1_3_0_65_sva_1;
  wire [3:0] s_output_1_19_16_46_sva_1;
  wire [3:0] s_output_1_19_16_31_sva_1;
  wire [3:0] s_output_1_3_0_35_sva_1;
  wire [3:0] s_output_1_19_16_61_sva_1;
  wire [3:0] s_output_1_3_0_50_sva_1;
  wire [3:0] s_output_1_3_0_20_sva_1;
  wire [3:0] s_output_1_19_16_17_sva_1;
  wire [3:0] s_output_1_3_0_66_sva_1;
  wire [3:0] s_output_1_19_16_47_sva_1;
  wire [3:0] s_output_1_19_16_32_sva_1;
  wire [3:0] s_output_1_3_0_36_sva_1;
  wire [3:0] s_output_1_19_16_62_sva_1;
  wire [3:0] s_output_1_3_0_51_sva_1;
  wire [3:0] s_output_1_3_0_21_sva_1;
  wire [3:0] s_output_1_19_16_18_sva_1;
  wire [3:0] s_output_1_3_0_67_sva_1;
  wire [3:0] s_output_1_19_16_48_sva_1;
  wire [3:0] s_output_1_19_16_33_sva_1;
  wire [3:0] s_output_1_3_0_37_sva_1;
  wire [3:0] s_output_1_19_16_63_sva_1;
  wire [3:0] s_output_1_3_0_52_sva_1;
  wire [3:0] s_output_1_3_0_22_sva_1;
  wire [3:0] s_output_1_3_0_5_sva_1;
  wire [3:0] s_output_1_19_16_1_sva_1;
  wire [3:0] s_output_1_19_16_3_sva_1;
  wire [3:0] s_output_1_19_16_sva_1;
  wire [3:0] s_output_1_3_0_7_sva_1;
  wire [3:0] s_output_1_19_16_2_sva_1;
  wire [3:0] s_output_1_3_0_sva_1;
  wire [3:0] s_output_1_3_0_6_sva_1;

  wire[0:0] loop_DES_rounds_1_xor_32_nl;
  wire[0:0] loop_DES_rounds_2_xor_32_nl;
  wire[0:0] loop_DES_rounds_1_xor_31_nl;
  wire[0:0] loop_DES_rounds_2_xor_31_nl;
  wire[0:0] loop_DES_rounds_1_xor_30_nl;
  wire[0:0] loop_DES_rounds_2_xor_30_nl;
  wire[0:0] loop_DES_rounds_1_xor_29_nl;
  wire[0:0] loop_DES_rounds_2_xor_29_nl;
  wire[0:0] loop_DES_rounds_1_xor_28_nl;
  wire[0:0] loop_DES_rounds_2_xor_28_nl;
  wire[0:0] loop_DES_rounds_1_xor_27_nl;
  wire[0:0] loop_DES_rounds_2_xor_27_nl;
  wire[0:0] loop_DES_rounds_1_xor_26_nl;
  wire[0:0] loop_DES_rounds_2_xor_26_nl;
  wire[0:0] loop_DES_rounds_1_xor_25_nl;
  wire[0:0] loop_DES_rounds_2_xor_25_nl;
  wire[0:0] loop_DES_rounds_1_xor_24_nl;
  wire[0:0] loop_DES_rounds_2_xor_24_nl;
  wire[0:0] loop_DES_rounds_1_xor_23_nl;
  wire[0:0] loop_DES_rounds_2_xor_23_nl;
  wire[0:0] loop_DES_rounds_1_xor_22_nl;
  wire[0:0] loop_DES_rounds_2_xor_22_nl;
  wire[0:0] loop_DES_rounds_1_xor_21_nl;
  wire[0:0] loop_DES_rounds_2_xor_21_nl;
  wire[0:0] loop_DES_rounds_1_xor_20_nl;
  wire[0:0] loop_DES_rounds_2_xor_20_nl;
  wire[0:0] loop_DES_rounds_1_xor_19_nl;
  wire[0:0] loop_DES_rounds_2_xor_19_nl;
  wire[0:0] loop_DES_rounds_1_xor_18_nl;
  wire[0:0] loop_DES_rounds_2_xor_18_nl;
  wire[0:0] loop_DES_rounds_1_xor_17_nl;
  wire[0:0] loop_DES_rounds_2_xor_17_nl;
  wire[0:0] loop_DES_rounds_1_xor_16_nl;
  wire[0:0] loop_DES_rounds_2_xor_16_nl;
  wire[0:0] loop_DES_rounds_1_xor_15_nl;
  wire[0:0] loop_DES_rounds_2_xor_15_nl;
  wire[0:0] loop_DES_rounds_1_xor_14_nl;
  wire[0:0] loop_DES_rounds_2_xor_14_nl;
  wire[0:0] loop_DES_rounds_1_xor_13_nl;
  wire[0:0] loop_DES_rounds_2_xor_13_nl;
  wire[0:0] loop_DES_rounds_1_xor_12_nl;
  wire[0:0] loop_DES_rounds_2_xor_12_nl;
  wire[0:0] loop_DES_rounds_1_xor_11_nl;
  wire[0:0] loop_DES_rounds_2_xor_11_nl;
  wire[0:0] loop_DES_rounds_1_xor_10_nl;
  wire[0:0] loop_DES_rounds_2_xor_10_nl;
  wire[0:0] loop_DES_rounds_1_xor_9_nl;
  wire[0:0] loop_DES_rounds_2_xor_9_nl;
  wire[0:0] loop_DES_rounds_1_xor_8_nl;
  wire[0:0] loop_DES_rounds_2_xor_8_nl;
  wire[0:0] loop_DES_rounds_1_xor_7_nl;
  wire[0:0] loop_DES_rounds_2_xor_7_nl;
  wire[0:0] loop_DES_rounds_1_xor_6_nl;
  wire[0:0] loop_DES_rounds_2_xor_6_nl;
  wire[0:0] loop_DES_rounds_1_xor_5_nl;
  wire[0:0] loop_DES_rounds_2_xor_5_nl;
  wire[0:0] loop_DES_rounds_1_xor_4_nl;
  wire[0:0] loop_DES_rounds_2_xor_4_nl;
  wire[0:0] loop_DES_rounds_1_xor_3_nl;
  wire[0:0] loop_DES_rounds_2_xor_3_nl;
  wire[0:0] loop_DES_rounds_1_xor_2_nl;
  wire[0:0] loop_DES_rounds_2_xor_2_nl;
  wire[0:0] loop_DES_rounds_1_xor_1_nl;
  wire[0:0] loop_DES_rounds_2_xor_1_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [63:0] nl_return_rsci_idat;
  assign nl_return_rsci_idat = {return_rsci_idat_63 , return_rsci_idat_62 , return_rsci_idat_61
      , return_rsci_idat_60 , return_rsci_idat_59 , return_rsci_idat_58 , return_rsci_idat_57
      , return_rsci_idat_56 , return_rsci_idat_55 , return_rsci_idat_54 , return_rsci_idat_53
      , return_rsci_idat_52 , return_rsci_idat_51 , return_rsci_idat_50 , return_rsci_idat_49
      , return_rsci_idat_48 , return_rsci_idat_47 , return_rsci_idat_46 , return_rsci_idat_45
      , return_rsci_idat_44 , return_rsci_idat_43 , return_rsci_idat_42 , return_rsci_idat_41
      , return_rsci_idat_40 , return_rsci_idat_39 , return_rsci_idat_38 , return_rsci_idat_37
      , return_rsci_idat_36 , return_rsci_idat_35 , return_rsci_idat_34 , return_rsci_idat_33
      , return_rsci_idat_32 , return_rsci_idat_31 , return_rsci_idat_30 , return_rsci_idat_29
      , return_rsci_idat_28 , return_rsci_idat_27 , return_rsci_idat_26 , return_rsci_idat_25
      , return_rsci_idat_24 , return_rsci_idat_23 , return_rsci_idat_22 , return_rsci_idat_21
      , return_rsci_idat_20 , return_rsci_idat_19 , return_rsci_idat_18 , return_rsci_idat_17
      , return_rsci_idat_16 , return_rsci_idat_15 , return_rsci_idat_14 , return_rsci_idat_13
      , return_rsci_idat_12 , return_rsci_idat_11 , return_rsci_idat_10 , return_rsci_idat_9
      , return_rsci_idat_8 , return_rsci_idat_7 , return_rsci_idat_6 , return_rsci_idat_5
      , return_rsci_idat_4 , return_rsci_idat_3 , return_rsci_idat_2 , return_rsci_idat_1
      , return_rsci_idat_0};
  wire[0:0] loop_DES_rounds_1_xor_50_nl;
  wire[0:0] loop_DES_rounds_1_xor_55_nl;
  wire[0:0] loop_DES_rounds_1_xor_51_nl;
  wire[0:0] loop_DES_rounds_1_xor_52_nl;
  wire[0:0] loop_DES_rounds_1_xor_53_nl;
  wire[0:0] loop_DES_rounds_1_xor_54_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_6_rg_addr;
  assign loop_DES_rounds_1_xor_50_nl = (input_rsci_idat[29]) ^ (key_rsci_idat[5]);
  assign loop_DES_rounds_1_xor_55_nl = (input_rsci_idat[3]) ^ (key_rsci_idat[23]);
  assign loop_DES_rounds_1_xor_51_nl = (input_rsci_idat[37]) ^ (key_rsci_idat[63]);
  assign loop_DES_rounds_1_xor_52_nl = (input_rsci_idat[45]) ^ (key_rsci_idat[28]);
  assign loop_DES_rounds_1_xor_53_nl = (input_rsci_idat[53]) ^ (key_rsci_idat[37]);
  assign loop_DES_rounds_1_xor_54_nl = (input_rsci_idat[61]) ^ (key_rsci_idat[46]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_6_rg_addr = {3'b011 , loop_DES_rounds_1_xor_50_nl
      , loop_DES_rounds_1_xor_55_nl , loop_DES_rounds_1_xor_51_nl , loop_DES_rounds_1_xor_52_nl
      , loop_DES_rounds_1_xor_53_nl , loop_DES_rounds_1_xor_54_nl};
  wire[0:0] loop_DES_rounds_1_xor_68_nl;
  wire[0:0] loop_DES_rounds_1_xor_73_nl;
  wire[0:0] loop_DES_rounds_1_xor_69_nl;
  wire[0:0] loop_DES_rounds_1_xor_70_nl;
  wire[0:0] loop_DES_rounds_1_xor_71_nl;
  wire[0:0] loop_DES_rounds_1_xor_72_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_5_rg_addr;
  assign loop_DES_rounds_1_xor_68_nl = (input_rsci_idat[59]) ^ (key_rsci_idat[3]);
  assign loop_DES_rounds_1_xor_73_nl = (input_rsci_idat[33]) ^ (key_rsci_idat[44]);
  assign loop_DES_rounds_1_xor_69_nl = (input_rsci_idat[1]) ^ (key_rsci_idat[43]);
  assign loop_DES_rounds_1_xor_70_nl = (input_rsci_idat[9]) ^ (key_rsci_idat[26]);
  assign loop_DES_rounds_1_xor_71_nl = (input_rsci_idat[17]) ^ (key_rsci_idat[1]);
  assign loop_DES_rounds_1_xor_72_nl = (input_rsci_idat[25]) ^ (key_rsci_idat[49]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_5_rg_addr = {3'b110 , loop_DES_rounds_1_xor_68_nl
      , loop_DES_rounds_1_xor_73_nl , loop_DES_rounds_1_xor_69_nl , loop_DES_rounds_1_xor_70_nl
      , loop_DES_rounds_1_xor_71_nl , loop_DES_rounds_1_xor_72_nl};
  wire[0:0] loop_DES_rounds_1_xor_38_nl;
  wire[0:0] loop_DES_rounds_1_xor_43_nl;
  wire[0:0] loop_DES_rounds_1_xor_39_nl;
  wire[0:0] loop_DES_rounds_1_xor_40_nl;
  wire[0:0] loop_DES_rounds_1_xor_41_nl;
  wire[0:0] loop_DES_rounds_1_xor_42_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_2_rg_addr;
  assign loop_DES_rounds_1_xor_38_nl = (input_rsci_idat[31]) ^ (key_rsci_idat[31]);
  assign loop_DES_rounds_1_xor_43_nl = (input_rsci_idat[5]) ^ (key_rsci_idat[22]);
  assign loop_DES_rounds_1_xor_39_nl = (input_rsci_idat[39]) ^ (key_rsci_idat[7]);
  assign loop_DES_rounds_1_xor_40_nl = (input_rsci_idat[47]) ^ (key_rsci_idat[62]);
  assign loop_DES_rounds_1_xor_41_nl = (input_rsci_idat[55]) ^ (key_rsci_idat[55]);
  assign loop_DES_rounds_1_xor_42_nl = (input_rsci_idat[63]) ^ (key_rsci_idat[45]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_2_rg_addr = {3'b001 , loop_DES_rounds_1_xor_38_nl
      , loop_DES_rounds_1_xor_43_nl , loop_DES_rounds_1_xor_39_nl , loop_DES_rounds_1_xor_40_nl
      , loop_DES_rounds_1_xor_41_nl , loop_DES_rounds_1_xor_42_nl};
  wire[0:0] loop_DES_rounds_1_xor_nl;
  wire[0:0] loop_DES_rounds_1_xor_37_nl;
  wire[0:0] loop_DES_rounds_1_xor_33_nl;
  wire[0:0] loop_DES_rounds_1_xor_34_nl;
  wire[0:0] loop_DES_rounds_1_xor_35_nl;
  wire[0:0] loop_DES_rounds_1_xor_36_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_rg_addr;
  assign loop_DES_rounds_1_xor_nl = (input_rsci_idat[57]) ^ (key_rsci_idat[54]);
  assign loop_DES_rounds_1_xor_37_nl = (input_rsci_idat[39]) ^ (key_rsci_idat[47]);
  assign loop_DES_rounds_1_xor_33_nl = (input_rsci_idat[7]) ^ (key_rsci_idat[13]);
  assign loop_DES_rounds_1_xor_34_nl = (input_rsci_idat[15]) ^ (key_rsci_idat[30]);
  assign loop_DES_rounds_1_xor_35_nl = (input_rsci_idat[23]) ^ (key_rsci_idat[4]);
  assign loop_DES_rounds_1_xor_36_nl = (input_rsci_idat[31]) ^ (key_rsci_idat[15]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_rg_addr = {3'b000 , loop_DES_rounds_1_xor_nl
      , loop_DES_rounds_1_xor_37_nl , loop_DES_rounds_1_xor_33_nl , loop_DES_rounds_1_xor_34_nl
      , loop_DES_rounds_1_xor_35_nl , loop_DES_rounds_1_xor_36_nl};
  wire[0:0] loop_DES_rounds_1_xor_56_nl;
  wire[0:0] loop_DES_rounds_1_xor_61_nl;
  wire[0:0] loop_DES_rounds_1_xor_57_nl;
  wire[0:0] loop_DES_rounds_1_xor_58_nl;
  wire[0:0] loop_DES_rounds_1_xor_59_nl;
  wire[0:0] loop_DES_rounds_1_xor_60_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_1_rg_addr;
  assign loop_DES_rounds_1_xor_56_nl = (input_rsci_idat[61]) ^ (key_rsci_idat[42]);
  assign loop_DES_rounds_1_xor_61_nl = (input_rsci_idat[35]) ^ (key_rsci_idat[60]);
  assign loop_DES_rounds_1_xor_57_nl = (input_rsci_idat[3]) ^ (key_rsci_idat[36]);
  assign loop_DES_rounds_1_xor_58_nl = (input_rsci_idat[11]) ^ (key_rsci_idat[25]);
  assign loop_DES_rounds_1_xor_59_nl = (input_rsci_idat[19]) ^ (key_rsci_idat[10]);
  assign loop_DES_rounds_1_xor_60_nl = (input_rsci_idat[27]) ^ (key_rsci_idat[27]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_1_rg_addr = {3'b100 , loop_DES_rounds_1_xor_56_nl
      , loop_DES_rounds_1_xor_61_nl , loop_DES_rounds_1_xor_57_nl , loop_DES_rounds_1_xor_58_nl
      , loop_DES_rounds_1_xor_59_nl , loop_DES_rounds_1_xor_60_nl};
  wire[0:0] loop_DES_rounds_1_xor_44_nl;
  wire[0:0] loop_DES_rounds_1_xor_49_nl;
  wire[0:0] loop_DES_rounds_1_xor_45_nl;
  wire[0:0] loop_DES_rounds_1_xor_46_nl;
  wire[0:0] loop_DES_rounds_1_xor_47_nl;
  wire[0:0] loop_DES_rounds_1_xor_48_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_4_rg_addr;
  assign loop_DES_rounds_1_xor_44_nl = (input_rsci_idat[63]) ^ (key_rsci_idat[61]);
  assign loop_DES_rounds_1_xor_49_nl = (input_rsci_idat[37]) ^ (key_rsci_idat[6]);
  assign loop_DES_rounds_1_xor_45_nl = (input_rsci_idat[5]) ^ (key_rsci_idat[29]);
  assign loop_DES_rounds_1_xor_46_nl = (input_rsci_idat[13]) ^ (key_rsci_idat[38]);
  assign loop_DES_rounds_1_xor_47_nl = (input_rsci_idat[21]) ^ (key_rsci_idat[39]);
  assign loop_DES_rounds_1_xor_48_nl = (input_rsci_idat[29]) ^ (key_rsci_idat[20]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_4_rg_addr = {3'b010 , loop_DES_rounds_1_xor_44_nl
      , loop_DES_rounds_1_xor_49_nl , loop_DES_rounds_1_xor_45_nl , loop_DES_rounds_1_xor_46_nl
      , loop_DES_rounds_1_xor_47_nl , loop_DES_rounds_1_xor_48_nl};
  wire[0:0] loop_DES_rounds_1_xor_62_nl;
  wire[0:0] loop_DES_rounds_1_xor_67_nl;
  wire[0:0] loop_DES_rounds_1_xor_63_nl;
  wire[0:0] loop_DES_rounds_1_xor_64_nl;
  wire[0:0] loop_DES_rounds_1_xor_65_nl;
  wire[0:0] loop_DES_rounds_1_xor_66_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_3_rg_addr;
  assign loop_DES_rounds_1_xor_62_nl = (input_rsci_idat[27]) ^ (key_rsci_idat[17]);
  assign loop_DES_rounds_1_xor_67_nl = (input_rsci_idat[1]) ^ (key_rsci_idat[35]);
  assign loop_DES_rounds_1_xor_63_nl = (input_rsci_idat[35]) ^ (key_rsci_idat[34]);
  assign loop_DES_rounds_1_xor_64_nl = (input_rsci_idat[43]) ^ (key_rsci_idat[59]);
  assign loop_DES_rounds_1_xor_65_nl = (input_rsci_idat[51]) ^ (key_rsci_idat[11]);
  assign loop_DES_rounds_1_xor_66_nl = (input_rsci_idat[59]) ^ (key_rsci_idat[41]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_3_rg_addr = {3'b101 , loop_DES_rounds_1_xor_62_nl
      , loop_DES_rounds_1_xor_67_nl , loop_DES_rounds_1_xor_63_nl , loop_DES_rounds_1_xor_64_nl
      , loop_DES_rounds_1_xor_65_nl , loop_DES_rounds_1_xor_66_nl};
  wire[0:0] loop_DES_rounds_1_xor_74_nl;
  wire[0:0] loop_DES_rounds_1_xor_79_nl;
  wire[0:0] loop_DES_rounds_1_xor_75_nl;
  wire[0:0] loop_DES_rounds_1_xor_76_nl;
  wire[0:0] loop_DES_rounds_1_xor_77_nl;
  wire[0:0] loop_DES_rounds_1_xor_78_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_7_rg_addr;
  assign loop_DES_rounds_1_xor_74_nl = (input_rsci_idat[25]) ^ (key_rsci_idat[19]);
  assign loop_DES_rounds_1_xor_79_nl = (input_rsci_idat[7]) ^ (key_rsci_idat[33]);
  assign loop_DES_rounds_1_xor_75_nl = (input_rsci_idat[33]) ^ (key_rsci_idat[50]);
  assign loop_DES_rounds_1_xor_76_nl = (input_rsci_idat[41]) ^ (key_rsci_idat[51]);
  assign loop_DES_rounds_1_xor_77_nl = (input_rsci_idat[49]) ^ (key_rsci_idat[2]);
  assign loop_DES_rounds_1_xor_78_nl = (input_rsci_idat[57]) ^ (key_rsci_idat[9]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_7_rg_addr = {3'b111 , loop_DES_rounds_1_xor_74_nl
      , loop_DES_rounds_1_xor_79_nl , loop_DES_rounds_1_xor_75_nl , loop_DES_rounds_1_xor_76_nl
      , loop_DES_rounds_1_xor_77_nl , loop_DES_rounds_1_xor_78_nl};
  wire[0:0] loop_DES_rounds_xor_nl;
  wire[0:0] loop_DES_rounds_xor_1_nl;
  wire[0:0] loop_DES_rounds_xor_2_nl;
  wire[0:0] loop_DES_rounds_xor_3_nl;
  wire[0:0] loop_DES_rounds_xor_4_nl;
  wire[0:0] loop_DES_rounds_xor_5_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_14_rg_addr;
  assign loop_DES_rounds_xor_nl = (input_sva[28]) ^ (s_output_1_3_0_53_sva[2]) ^
      (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_xor_1_nl = (input_sva[2]) ^ (s_output_1_19_16_19_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign loop_DES_rounds_xor_2_nl = (input_sva[36]) ^ (s_output_1_19_16_34_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_xor_3_nl = (input_sva[44]) ^ (s_output_1_3_0_23_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_xor_4_nl = (input_sva[52]) ^ (s_output_1_3_0_8_sva[1]) ^
      (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_xor_5_nl = (input_sva[60]) ^ (s_output_1_19_16_49_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_14_rg_addr = {3'b011 , loop_DES_rounds_xor_nl
      , loop_DES_rounds_xor_1_nl , loop_DES_rounds_xor_2_nl , loop_DES_rounds_xor_3_nl
      , loop_DES_rounds_xor_4_nl , loop_DES_rounds_xor_5_nl};
  wire[0:0] loop_DES_rounds_xor_6_nl;
  wire[0:0] loop_DES_rounds_xor_7_nl;
  wire[0:0] loop_DES_rounds_xor_8_nl;
  wire[0:0] loop_DES_rounds_xor_9_nl;
  wire[0:0] loop_DES_rounds_xor_10_nl;
  wire[0:0] loop_DES_rounds_xor_11_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_13_rg_addr;
  assign loop_DES_rounds_xor_6_nl = (input_sva[58]) ^ (s_output_1_19_16_49_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_xor_7_nl = (input_sva[32]) ^ (s_output_1_3_0_38_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_xor_8_nl = (input_sva[0]) ^ (s_output_1_3_0_23_sva[1]) ^
      (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_xor_9_nl = (input_sva[8]) ^ (s_output_1_19_16_4_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_xor_10_nl = (input_sva[16]) ^ (s_output_1_3_0_8_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_xor_11_nl = (input_sva[24]) ^ (s_output_1_19_16_34_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_13_rg_addr = {3'b110 , loop_DES_rounds_xor_6_nl
      , loop_DES_rounds_xor_7_nl , loop_DES_rounds_xor_8_nl , loop_DES_rounds_xor_9_nl
      , loop_DES_rounds_xor_10_nl , loop_DES_rounds_xor_11_nl};
  wire[0:0] loop_DES_rounds_xor_12_nl;
  wire[0:0] loop_DES_rounds_xor_13_nl;
  wire[0:0] loop_DES_rounds_xor_14_nl;
  wire[0:0] loop_DES_rounds_xor_15_nl;
  wire[0:0] loop_DES_rounds_xor_16_nl;
  wire[0:0] loop_DES_rounds_xor_17_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_10_rg_addr;
  assign loop_DES_rounds_xor_12_nl = (input_sva[30]) ^ (s_output_1_3_0_38_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_xor_13_nl = (input_sva[4]) ^ (s_output_1_19_16_19_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_xor_14_nl = (input_sva[38]) ^ (s_output_1_3_0_8_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign loop_DES_rounds_xor_15_nl = (input_sva[46]) ^ (s_output_1_19_16_49_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign loop_DES_rounds_xor_16_nl = (input_sva[54]) ^ (s_output_1_3_0_53_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_xor_17_nl = (input_sva[62]) ^ (s_output_1_3_0_23_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_10_rg_addr = {3'b001 , loop_DES_rounds_xor_12_nl
      , loop_DES_rounds_xor_13_nl , loop_DES_rounds_xor_14_nl , loop_DES_rounds_xor_15_nl
      , loop_DES_rounds_xor_16_nl , loop_DES_rounds_xor_17_nl};
  wire[0:0] loop_DES_rounds_xor_18_nl;
  wire[0:0] loop_DES_rounds_xor_19_nl;
  wire[0:0] loop_DES_rounds_xor_20_nl;
  wire[0:0] loop_DES_rounds_xor_21_nl;
  wire[0:0] loop_DES_rounds_xor_22_nl;
  wire[0:0] loop_DES_rounds_xor_23_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_8_rg_addr;
  assign loop_DES_rounds_xor_18_nl = (input_sva[56]) ^ (s_output_1_3_0_53_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_xor_19_nl = (input_sva[38]) ^ (s_output_1_3_0_8_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_xor_20_nl = (input_sva[6]) ^ (s_output_1_19_16_4_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_xor_21_nl = (input_sva[14]) ^ (s_output_1_19_16_34_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign loop_DES_rounds_xor_22_nl = (input_sva[22]) ^ (s_output_1_3_0_23_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_xor_23_nl = (input_sva[30]) ^ (s_output_1_3_0_38_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_8_rg_addr = {3'b000 , loop_DES_rounds_xor_18_nl
      , loop_DES_rounds_xor_19_nl , loop_DES_rounds_xor_20_nl , loop_DES_rounds_xor_21_nl
      , loop_DES_rounds_xor_22_nl , loop_DES_rounds_xor_23_nl};
  wire[0:0] loop_DES_rounds_xor_24_nl;
  wire[0:0] loop_DES_rounds_xor_25_nl;
  wire[0:0] loop_DES_rounds_xor_26_nl;
  wire[0:0] loop_DES_rounds_xor_27_nl;
  wire[0:0] loop_DES_rounds_xor_28_nl;
  wire[0:0] loop_DES_rounds_xor_29_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_9_rg_addr;
  assign loop_DES_rounds_xor_24_nl = (input_sva[60]) ^ (s_output_1_19_16_49_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_xor_25_nl = (input_sva[34]) ^ (s_output_1_3_0_8_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_xor_26_nl = (input_sva[2]) ^ (s_output_1_19_16_19_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_xor_27_nl = (input_sva[10]) ^ (s_output_1_19_16_34_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_xor_28_nl = (input_sva[18]) ^ (s_output_1_3_0_38_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_xor_29_nl = (input_sva[26]) ^ (s_output_1_19_16_4_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_9_rg_addr = {3'b100 , loop_DES_rounds_xor_24_nl
      , loop_DES_rounds_xor_25_nl , loop_DES_rounds_xor_26_nl , loop_DES_rounds_xor_27_nl
      , loop_DES_rounds_xor_28_nl , loop_DES_rounds_xor_29_nl};
  wire[0:0] loop_DES_rounds_xor_30_nl;
  wire[0:0] loop_DES_rounds_xor_31_nl;
  wire[0:0] loop_DES_rounds_xor_32_nl;
  wire[0:0] loop_DES_rounds_xor_33_nl;
  wire[0:0] loop_DES_rounds_xor_34_nl;
  wire[0:0] loop_DES_rounds_xor_35_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_12_rg_addr;
  assign loop_DES_rounds_xor_30_nl = (input_sva[62]) ^ (s_output_1_3_0_23_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_xor_31_nl = (input_sva[36]) ^ (s_output_1_19_16_34_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_xor_32_nl = (input_sva[4]) ^ (s_output_1_19_16_19_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_xor_33_nl = (input_sva[12]) ^ (s_output_1_19_16_4_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_xor_34_nl = (input_sva[20]) ^ (s_output_1_3_0_38_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_xor_35_nl = (input_sva[28]) ^ (s_output_1_3_0_53_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_12_rg_addr = {3'b010 , loop_DES_rounds_xor_30_nl
      , loop_DES_rounds_xor_31_nl , loop_DES_rounds_xor_32_nl , loop_DES_rounds_xor_33_nl
      , loop_DES_rounds_xor_34_nl , loop_DES_rounds_xor_35_nl};
  wire[0:0] loop_DES_rounds_xor_36_nl;
  wire[0:0] loop_DES_rounds_xor_37_nl;
  wire[0:0] loop_DES_rounds_xor_38_nl;
  wire[0:0] loop_DES_rounds_xor_39_nl;
  wire[0:0] loop_DES_rounds_xor_40_nl;
  wire[0:0] loop_DES_rounds_xor_41_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_11_rg_addr;
  assign loop_DES_rounds_xor_36_nl = (input_sva[26]) ^ (s_output_1_19_16_4_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_xor_37_nl = (input_sva[0]) ^ (s_output_1_3_0_23_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_xor_38_nl = (key_io_read_key_rsc_cse_63_1_sva[41]) ^ (input_sva[34])
      ^ (s_output_1_3_0_8_sva[0]);
  assign loop_DES_rounds_xor_39_nl = (input_sva[42]) ^ (s_output_1_3_0_53_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_xor_40_nl = (input_sva[50]) ^ (s_output_1_19_16_19_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_xor_41_nl = (input_sva[58]) ^ (s_output_1_19_16_49_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_11_rg_addr = {3'b101 , loop_DES_rounds_xor_36_nl
      , loop_DES_rounds_xor_37_nl , loop_DES_rounds_xor_38_nl , loop_DES_rounds_xor_39_nl
      , loop_DES_rounds_xor_40_nl , loop_DES_rounds_xor_41_nl};
  wire[0:0] loop_DES_rounds_xor_42_nl;
  wire[0:0] loop_DES_rounds_xor_43_nl;
  wire[0:0] loop_DES_rounds_xor_44_nl;
  wire[0:0] loop_DES_rounds_xor_45_nl;
  wire[0:0] loop_DES_rounds_xor_46_nl;
  wire[0:0] loop_DES_rounds_xor_47_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_15_rg_addr;
  assign loop_DES_rounds_xor_42_nl = (input_sva[24]) ^ (s_output_1_19_16_34_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_xor_43_nl = (input_sva[6]) ^ (s_output_1_19_16_4_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_xor_44_nl = (input_sva[32]) ^ (s_output_1_3_0_38_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_xor_45_nl = (input_sva[40]) ^ (s_output_1_19_16_49_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_xor_46_nl = (input_sva[48]) ^ (s_output_1_19_16_19_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_xor_47_nl = (input_sva[56]) ^ (s_output_1_3_0_53_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_15_rg_addr = {3'b111 , loop_DES_rounds_xor_42_nl
      , loop_DES_rounds_xor_43_nl , loop_DES_rounds_xor_44_nl , loop_DES_rounds_xor_45_nl
      , loop_DES_rounds_xor_46_nl , loop_DES_rounds_xor_47_nl};
  wire[0:0] loop_DES_rounds_xor_48_nl;
  wire[0:0] loop_DES_rounds_xor_49_nl;
  wire[0:0] loop_DES_rounds_xor_50_nl;
  wire[0:0] loop_DES_rounds_xor_51_nl;
  wire[0:0] loop_DES_rounds_xor_52_nl;
  wire[0:0] loop_DES_rounds_xor_53_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_22_rg_addr;
  assign loop_DES_rounds_xor_48_nl = (key_io_read_key_rsc_cse_63_1_sva[28]) ^ (input_sva[29])
      ^ (s_output_1_3_0_54_sva[2]);
  assign loop_DES_rounds_xor_49_nl = (input_sva[3]) ^ (s_output_1_19_16_20_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_xor_50_nl = (key_io_read_key_rsc_cse_63_1_sva[21]) ^ (input_sva[37])
      ^ (s_output_1_19_16_35_sva[3]);
  assign loop_DES_rounds_xor_51_nl = (input_sva[45]) ^ (s_output_1_3_0_24_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_xor_52_nl = (input_sva[53]) ^ (s_output_1_3_0_9_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_xor_53_nl = (input_sva[61]) ^ (s_output_1_19_16_50_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_22_rg_addr = {3'b011 , loop_DES_rounds_xor_48_nl
      , loop_DES_rounds_xor_49_nl , loop_DES_rounds_xor_50_nl , loop_DES_rounds_xor_51_nl
      , loop_DES_rounds_xor_52_nl , loop_DES_rounds_xor_53_nl};
  wire[0:0] loop_DES_rounds_xor_54_nl;
  wire[0:0] loop_DES_rounds_xor_55_nl;
  wire[0:0] loop_DES_rounds_xor_56_nl;
  wire[0:0] loop_DES_rounds_xor_57_nl;
  wire[0:0] loop_DES_rounds_xor_58_nl;
  wire[0:0] loop_DES_rounds_xor_59_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_21_rg_addr;
  assign loop_DES_rounds_xor_54_nl = (input_sva[59]) ^ (s_output_1_19_16_50_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_xor_55_nl = (input_sva[33]) ^ (s_output_1_3_0_39_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_xor_56_nl = (input_sva[1]) ^ (s_output_1_3_0_24_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_xor_57_nl = (input_sva[9]) ^ (s_output_1_19_16_5_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_xor_58_nl = (input_sva[17]) ^ (s_output_1_3_0_9_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_xor_59_nl = (input_sva[25]) ^ (s_output_1_19_16_35_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_21_rg_addr = {3'b110 , loop_DES_rounds_xor_54_nl
      , loop_DES_rounds_xor_55_nl , loop_DES_rounds_xor_56_nl , loop_DES_rounds_xor_57_nl
      , loop_DES_rounds_xor_58_nl , loop_DES_rounds_xor_59_nl};
  wire[0:0] loop_DES_rounds_xor_60_nl;
  wire[0:0] loop_DES_rounds_xor_61_nl;
  wire[0:0] loop_DES_rounds_xor_62_nl;
  wire[0:0] loop_DES_rounds_xor_63_nl;
  wire[0:0] loop_DES_rounds_xor_64_nl;
  wire[0:0] loop_DES_rounds_xor_65_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_18_rg_addr;
  assign loop_DES_rounds_xor_60_nl = (input_sva[31]) ^ (s_output_1_3_0_39_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_xor_61_nl = (input_sva[5]) ^ (s_output_1_19_16_20_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_xor_62_nl = (input_sva[39]) ^ (s_output_1_3_0_9_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign loop_DES_rounds_xor_63_nl = (input_sva[47]) ^ (s_output_1_19_16_50_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_xor_64_nl = (input_sva[55]) ^ (s_output_1_3_0_54_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_xor_65_nl = (input_sva[63]) ^ (s_output_1_3_0_24_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_18_rg_addr = {3'b001 , loop_DES_rounds_xor_60_nl
      , loop_DES_rounds_xor_61_nl , loop_DES_rounds_xor_62_nl , loop_DES_rounds_xor_63_nl
      , loop_DES_rounds_xor_64_nl , loop_DES_rounds_xor_65_nl};
  wire[0:0] loop_DES_rounds_xor_66_nl;
  wire[0:0] loop_DES_rounds_xor_67_nl;
  wire[0:0] loop_DES_rounds_xor_68_nl;
  wire[0:0] loop_DES_rounds_xor_69_nl;
  wire[0:0] loop_DES_rounds_xor_70_nl;
  wire[0:0] loop_DES_rounds_xor_71_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_16_rg_addr;
  assign loop_DES_rounds_xor_66_nl = (input_sva[57]) ^ (s_output_1_3_0_54_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_xor_67_nl = (input_sva[39]) ^ (s_output_1_3_0_9_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_xor_68_nl = (input_sva[7]) ^ (s_output_1_19_16_5_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_xor_69_nl = (input_sva[15]) ^ (s_output_1_19_16_35_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign loop_DES_rounds_xor_70_nl = (input_sva[23]) ^ (s_output_1_3_0_24_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign loop_DES_rounds_xor_71_nl = (input_sva[31]) ^ (s_output_1_3_0_39_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_16_rg_addr = {3'b000 , loop_DES_rounds_xor_66_nl
      , loop_DES_rounds_xor_67_nl , loop_DES_rounds_xor_68_nl , loop_DES_rounds_xor_69_nl
      , loop_DES_rounds_xor_70_nl , loop_DES_rounds_xor_71_nl};
  wire[0:0] loop_DES_rounds_xor_72_nl;
  wire[0:0] loop_DES_rounds_xor_73_nl;
  wire[0:0] loop_DES_rounds_xor_74_nl;
  wire[0:0] loop_DES_rounds_xor_75_nl;
  wire[0:0] loop_DES_rounds_xor_76_nl;
  wire[0:0] loop_DES_rounds_xor_77_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_17_rg_addr;
  assign loop_DES_rounds_xor_72_nl = (key_io_read_key_rsc_cse_63_1_sva[2]) ^ (input_sva[61])
      ^ (s_output_1_19_16_50_sva[2]);
  assign loop_DES_rounds_xor_73_nl = (input_sva[35]) ^ (s_output_1_3_0_9_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_xor_74_nl = (key_io_read_key_rsc_cse_63_1_sva[59]) ^ (input_sva[3])
      ^ (s_output_1_19_16_20_sva[2]);
  assign loop_DES_rounds_xor_75_nl = (input_sva[11]) ^ (s_output_1_19_16_35_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_xor_76_nl = (input_sva[19]) ^ (s_output_1_3_0_39_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_xor_77_nl = (input_sva[27]) ^ (s_output_1_19_16_5_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_17_rg_addr = {3'b100 , loop_DES_rounds_xor_72_nl
      , loop_DES_rounds_xor_73_nl , loop_DES_rounds_xor_74_nl , loop_DES_rounds_xor_75_nl
      , loop_DES_rounds_xor_76_nl , loop_DES_rounds_xor_77_nl};
  wire[0:0] loop_DES_rounds_xor_78_nl;
  wire[0:0] loop_DES_rounds_xor_79_nl;
  wire[0:0] loop_DES_rounds_xor_80_nl;
  wire[0:0] loop_DES_rounds_xor_81_nl;
  wire[0:0] loop_DES_rounds_xor_82_nl;
  wire[0:0] loop_DES_rounds_xor_83_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_20_rg_addr;
  assign loop_DES_rounds_xor_78_nl = (key_io_read_key_rsc_cse_63_1_sva[19]) ^ (input_sva[63])
      ^ (s_output_1_3_0_24_sva[3]);
  assign loop_DES_rounds_xor_79_nl = (input_sva[37]) ^ (s_output_1_19_16_35_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_xor_80_nl = (input_sva[5]) ^ (s_output_1_19_16_20_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_xor_81_nl = (input_sva[13]) ^ (s_output_1_19_16_5_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_xor_82_nl = (input_sva[21]) ^ (s_output_1_3_0_39_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_xor_83_nl = (input_sva[29]) ^ (s_output_1_3_0_54_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_20_rg_addr = {3'b010 , loop_DES_rounds_xor_78_nl
      , loop_DES_rounds_xor_79_nl , loop_DES_rounds_xor_80_nl , loop_DES_rounds_xor_81_nl
      , loop_DES_rounds_xor_82_nl , loop_DES_rounds_xor_83_nl};
  wire[0:0] loop_DES_rounds_xor_84_nl;
  wire[0:0] loop_DES_rounds_xor_85_nl;
  wire[0:0] loop_DES_rounds_xor_86_nl;
  wire[0:0] loop_DES_rounds_xor_87_nl;
  wire[0:0] loop_DES_rounds_xor_88_nl;
  wire[0:0] loop_DES_rounds_xor_89_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_19_rg_addr;
  assign loop_DES_rounds_xor_84_nl = (input_sva[27]) ^ (s_output_1_19_16_5_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_xor_85_nl = (input_sva[1]) ^ (s_output_1_3_0_24_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_xor_86_nl = (input_sva[35]) ^ (s_output_1_3_0_9_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_xor_87_nl = (input_sva[43]) ^ (s_output_1_3_0_54_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_xor_88_nl = (input_sva[51]) ^ (s_output_1_19_16_20_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_xor_89_nl = (key_io_read_key_rsc_cse_63_1_sva[1]) ^ (input_sva[59])
      ^ (s_output_1_19_16_50_sva[3]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_19_rg_addr = {3'b101 , loop_DES_rounds_xor_84_nl
      , loop_DES_rounds_xor_85_nl , loop_DES_rounds_xor_86_nl , loop_DES_rounds_xor_87_nl
      , loop_DES_rounds_xor_88_nl , loop_DES_rounds_xor_89_nl};
  wire[0:0] loop_DES_rounds_xor_90_nl;
  wire[0:0] loop_DES_rounds_xor_91_nl;
  wire[0:0] loop_DES_rounds_xor_92_nl;
  wire[0:0] loop_DES_rounds_xor_93_nl;
  wire[0:0] loop_DES_rounds_xor_94_nl;
  wire[0:0] loop_DES_rounds_xor_95_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_23_rg_addr;
  assign loop_DES_rounds_xor_90_nl = (input_sva[25]) ^ (s_output_1_19_16_35_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_xor_91_nl = (input_sva[7]) ^ (s_output_1_19_16_5_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign loop_DES_rounds_xor_92_nl = (input_sva[33]) ^ (s_output_1_3_0_39_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_xor_93_nl = (input_sva[41]) ^ (s_output_1_19_16_50_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_xor_94_nl = (input_sva[49]) ^ (s_output_1_19_16_20_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign loop_DES_rounds_xor_95_nl = (input_sva[57]) ^ (s_output_1_3_0_54_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_23_rg_addr = {3'b111 , loop_DES_rounds_xor_90_nl
      , loop_DES_rounds_xor_91_nl , loop_DES_rounds_xor_92_nl , loop_DES_rounds_xor_93_nl
      , loop_DES_rounds_xor_94_nl , loop_DES_rounds_xor_95_nl};
  wire[0:0] loop_DES_rounds_4_xor_50_nl;
  wire[0:0] loop_DES_rounds_4_xor_55_nl;
  wire[0:0] loop_DES_rounds_4_xor_51_nl;
  wire[0:0] loop_DES_rounds_4_xor_52_nl;
  wire[0:0] loop_DES_rounds_4_xor_53_nl;
  wire[0:0] loop_DES_rounds_4_xor_54_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_30_rg_addr;
  assign loop_DES_rounds_4_xor_50_nl = R_20_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_4_xor_55_nl = R_15_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_4_xor_51_nl = R_19_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign loop_DES_rounds_4_xor_52_nl = R_18_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_4_xor_53_nl = R_17_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_4_xor_54_nl = R_16_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_30_rg_addr = {3'b011 , loop_DES_rounds_4_xor_50_nl
      , loop_DES_rounds_4_xor_55_nl , loop_DES_rounds_4_xor_51_nl , loop_DES_rounds_4_xor_52_nl
      , loop_DES_rounds_4_xor_53_nl , loop_DES_rounds_4_xor_54_nl};
  wire[0:0] loop_DES_rounds_4_xor_68_nl;
  wire[0:0] loop_DES_rounds_4_xor_73_nl;
  wire[0:0] loop_DES_rounds_4_xor_69_nl;
  wire[0:0] loop_DES_rounds_4_xor_70_nl;
  wire[0:0] loop_DES_rounds_4_xor_71_nl;
  wire[0:0] loop_DES_rounds_4_xor_72_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_29_rg_addr;
  assign loop_DES_rounds_4_xor_68_nl = R_8_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_4_xor_73_nl = R_3_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_4_xor_69_nl = R_7_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_4_xor_70_nl = R_6_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_4_xor_71_nl = R_5_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_4_xor_72_nl = R_4_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_29_rg_addr = {3'b110 , loop_DES_rounds_4_xor_68_nl
      , loop_DES_rounds_4_xor_73_nl , loop_DES_rounds_4_xor_69_nl , loop_DES_rounds_4_xor_70_nl
      , loop_DES_rounds_4_xor_71_nl , loop_DES_rounds_4_xor_72_nl};
  wire[0:0] loop_DES_rounds_4_xor_38_nl;
  wire[0:0] loop_DES_rounds_4_xor_43_nl;
  wire[0:0] loop_DES_rounds_4_xor_39_nl;
  wire[0:0] loop_DES_rounds_4_xor_40_nl;
  wire[0:0] loop_DES_rounds_4_xor_41_nl;
  wire[0:0] loop_DES_rounds_4_xor_42_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_26_rg_addr;
  assign loop_DES_rounds_4_xor_38_nl = R_28_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_4_xor_43_nl = R_23_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_4_xor_39_nl = R_27_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_4_xor_40_nl = R_26_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_4_xor_41_nl = R_25_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_4_xor_42_nl = R_24_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_26_rg_addr = {3'b001 , loop_DES_rounds_4_xor_38_nl
      , loop_DES_rounds_4_xor_43_nl , loop_DES_rounds_4_xor_39_nl , loop_DES_rounds_4_xor_40_nl
      , loop_DES_rounds_4_xor_41_nl , loop_DES_rounds_4_xor_42_nl};
  wire[0:0] loop_DES_rounds_4_xor_nl;
  wire[0:0] loop_DES_rounds_4_xor_37_nl;
  wire[0:0] loop_DES_rounds_4_xor_33_nl;
  wire[0:0] loop_DES_rounds_4_xor_34_nl;
  wire[0:0] loop_DES_rounds_4_xor_35_nl;
  wire[0:0] loop_DES_rounds_4_xor_36_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_24_rg_addr;
  assign loop_DES_rounds_4_xor_nl = R_0_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign loop_DES_rounds_4_xor_37_nl = R_27_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign loop_DES_rounds_4_xor_33_nl = R_31_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_4_xor_34_nl = R_30_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign loop_DES_rounds_4_xor_35_nl = R_29_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign loop_DES_rounds_4_xor_36_nl = R_28_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_24_rg_addr = {3'b000 , loop_DES_rounds_4_xor_nl
      , loop_DES_rounds_4_xor_37_nl , loop_DES_rounds_4_xor_33_nl , loop_DES_rounds_4_xor_34_nl
      , loop_DES_rounds_4_xor_35_nl , loop_DES_rounds_4_xor_36_nl};
  wire[0:0] loop_DES_rounds_4_xor_56_nl;
  wire[0:0] loop_DES_rounds_4_xor_61_nl;
  wire[0:0] loop_DES_rounds_4_xor_57_nl;
  wire[0:0] loop_DES_rounds_4_xor_58_nl;
  wire[0:0] loop_DES_rounds_4_xor_59_nl;
  wire[0:0] loop_DES_rounds_4_xor_60_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_25_rg_addr;
  assign loop_DES_rounds_4_xor_56_nl = R_16_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_4_xor_61_nl = R_11_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_4_xor_57_nl = R_15_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_4_xor_58_nl = R_14_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_4_xor_59_nl = R_13_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_4_xor_60_nl = R_12_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_25_rg_addr = {3'b100 , loop_DES_rounds_4_xor_56_nl
      , loop_DES_rounds_4_xor_61_nl , loop_DES_rounds_4_xor_57_nl , loop_DES_rounds_4_xor_58_nl
      , loop_DES_rounds_4_xor_59_nl , loop_DES_rounds_4_xor_60_nl};
  wire[0:0] loop_DES_rounds_4_xor_44_nl;
  wire[0:0] loop_DES_rounds_4_xor_49_nl;
  wire[0:0] loop_DES_rounds_4_xor_45_nl;
  wire[0:0] loop_DES_rounds_4_xor_46_nl;
  wire[0:0] loop_DES_rounds_4_xor_47_nl;
  wire[0:0] loop_DES_rounds_4_xor_48_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_28_rg_addr;
  assign loop_DES_rounds_4_xor_44_nl = R_24_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_4_xor_49_nl = R_19_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_4_xor_45_nl = R_23_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_4_xor_46_nl = R_22_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_4_xor_47_nl = R_21_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_4_xor_48_nl = R_20_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_28_rg_addr = {3'b010 , loop_DES_rounds_4_xor_44_nl
      , loop_DES_rounds_4_xor_49_nl , loop_DES_rounds_4_xor_45_nl , loop_DES_rounds_4_xor_46_nl
      , loop_DES_rounds_4_xor_47_nl , loop_DES_rounds_4_xor_48_nl};
  wire[0:0] loop_DES_rounds_4_xor_62_nl;
  wire[0:0] loop_DES_rounds_4_xor_67_nl;
  wire[0:0] loop_DES_rounds_4_xor_63_nl;
  wire[0:0] loop_DES_rounds_4_xor_64_nl;
  wire[0:0] loop_DES_rounds_4_xor_65_nl;
  wire[0:0] loop_DES_rounds_4_xor_66_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_27_rg_addr;
  assign loop_DES_rounds_4_xor_62_nl = R_12_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign loop_DES_rounds_4_xor_67_nl = R_7_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_4_xor_63_nl = R_11_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_4_xor_64_nl = R_10_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_4_xor_65_nl = R_9_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_4_xor_66_nl = R_8_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_27_rg_addr = {3'b101 , loop_DES_rounds_4_xor_62_nl
      , loop_DES_rounds_4_xor_67_nl , loop_DES_rounds_4_xor_63_nl , loop_DES_rounds_4_xor_64_nl
      , loop_DES_rounds_4_xor_65_nl , loop_DES_rounds_4_xor_66_nl};
  wire[0:0] loop_DES_rounds_4_xor_74_nl;
  wire[0:0] loop_DES_rounds_4_xor_79_nl;
  wire[0:0] loop_DES_rounds_4_xor_75_nl;
  wire[0:0] loop_DES_rounds_4_xor_76_nl;
  wire[0:0] loop_DES_rounds_4_xor_77_nl;
  wire[0:0] loop_DES_rounds_4_xor_78_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_31_rg_addr;
  assign loop_DES_rounds_4_xor_74_nl = R_4_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_4_xor_79_nl = R_31_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_4_xor_75_nl = R_3_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_4_xor_76_nl = R_2_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_4_xor_77_nl = R_1_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_4_xor_78_nl = R_0_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_31_rg_addr = {3'b111 , loop_DES_rounds_4_xor_74_nl
      , loop_DES_rounds_4_xor_79_nl , loop_DES_rounds_4_xor_75_nl , loop_DES_rounds_4_xor_76_nl
      , loop_DES_rounds_4_xor_77_nl , loop_DES_rounds_4_xor_78_nl};
  wire[0:0] loop_DES_rounds_5_xor_50_nl;
  wire[0:0] loop_DES_rounds_5_xor_55_nl;
  wire[0:0] loop_DES_rounds_5_xor_51_nl;
  wire[0:0] loop_DES_rounds_5_xor_52_nl;
  wire[0:0] loop_DES_rounds_5_xor_53_nl;
  wire[0:0] loop_DES_rounds_5_xor_54_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_38_rg_addr;
  assign loop_DES_rounds_5_xor_50_nl = R_20_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_5_xor_55_nl = R_15_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_5_xor_51_nl = R_19_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign loop_DES_rounds_5_xor_52_nl = R_18_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_5_xor_53_nl = R_17_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign loop_DES_rounds_5_xor_54_nl = R_16_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_38_rg_addr = {3'b011 , loop_DES_rounds_5_xor_50_nl
      , loop_DES_rounds_5_xor_55_nl , loop_DES_rounds_5_xor_51_nl , loop_DES_rounds_5_xor_52_nl
      , loop_DES_rounds_5_xor_53_nl , loop_DES_rounds_5_xor_54_nl};
  wire[0:0] loop_DES_rounds_5_xor_68_nl;
  wire[0:0] loop_DES_rounds_5_xor_73_nl;
  wire[0:0] loop_DES_rounds_5_xor_69_nl;
  wire[0:0] loop_DES_rounds_5_xor_70_nl;
  wire[0:0] loop_DES_rounds_5_xor_71_nl;
  wire[0:0] loop_DES_rounds_5_xor_72_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_37_rg_addr;
  assign loop_DES_rounds_5_xor_68_nl = R_8_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_5_xor_73_nl = R_3_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_5_xor_69_nl = R_7_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_5_xor_70_nl = R_6_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_5_xor_71_nl = R_5_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign loop_DES_rounds_5_xor_72_nl = R_4_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_37_rg_addr = {3'b110 , loop_DES_rounds_5_xor_68_nl
      , loop_DES_rounds_5_xor_73_nl , loop_DES_rounds_5_xor_69_nl , loop_DES_rounds_5_xor_70_nl
      , loop_DES_rounds_5_xor_71_nl , loop_DES_rounds_5_xor_72_nl};
  wire[0:0] loop_DES_rounds_5_xor_38_nl;
  wire[0:0] loop_DES_rounds_5_xor_43_nl;
  wire[0:0] loop_DES_rounds_5_xor_39_nl;
  wire[0:0] loop_DES_rounds_5_xor_40_nl;
  wire[0:0] loop_DES_rounds_5_xor_41_nl;
  wire[0:0] loop_DES_rounds_5_xor_42_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_34_rg_addr;
  assign loop_DES_rounds_5_xor_38_nl = R_28_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign loop_DES_rounds_5_xor_43_nl = R_23_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_5_xor_39_nl = R_27_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_5_xor_40_nl = R_26_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_5_xor_41_nl = R_25_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_5_xor_42_nl = R_24_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_34_rg_addr = {3'b001 , loop_DES_rounds_5_xor_38_nl
      , loop_DES_rounds_5_xor_43_nl , loop_DES_rounds_5_xor_39_nl , loop_DES_rounds_5_xor_40_nl
      , loop_DES_rounds_5_xor_41_nl , loop_DES_rounds_5_xor_42_nl};
  wire[0:0] loop_DES_rounds_5_xor_nl;
  wire[0:0] loop_DES_rounds_5_xor_37_nl;
  wire[0:0] loop_DES_rounds_5_xor_33_nl;
  wire[0:0] loop_DES_rounds_5_xor_34_nl;
  wire[0:0] loop_DES_rounds_5_xor_35_nl;
  wire[0:0] loop_DES_rounds_5_xor_36_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_32_rg_addr;
  assign loop_DES_rounds_5_xor_nl = R_0_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_5_xor_37_nl = R_27_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign loop_DES_rounds_5_xor_33_nl = R_31_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_5_xor_34_nl = R_30_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_5_xor_35_nl = R_29_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign loop_DES_rounds_5_xor_36_nl = R_28_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_32_rg_addr = {3'b000 , loop_DES_rounds_5_xor_nl
      , loop_DES_rounds_5_xor_37_nl , loop_DES_rounds_5_xor_33_nl , loop_DES_rounds_5_xor_34_nl
      , loop_DES_rounds_5_xor_35_nl , loop_DES_rounds_5_xor_36_nl};
  wire[0:0] loop_DES_rounds_5_xor_56_nl;
  wire[0:0] loop_DES_rounds_5_xor_61_nl;
  wire[0:0] loop_DES_rounds_5_xor_57_nl;
  wire[0:0] loop_DES_rounds_5_xor_58_nl;
  wire[0:0] loop_DES_rounds_5_xor_59_nl;
  wire[0:0] loop_DES_rounds_5_xor_60_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_33_rg_addr;
  assign loop_DES_rounds_5_xor_56_nl = R_16_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_5_xor_61_nl = R_11_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_5_xor_57_nl = R_15_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_5_xor_58_nl = R_14_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_5_xor_59_nl = R_13_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_5_xor_60_nl = R_12_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_33_rg_addr = {3'b100 , loop_DES_rounds_5_xor_56_nl
      , loop_DES_rounds_5_xor_61_nl , loop_DES_rounds_5_xor_57_nl , loop_DES_rounds_5_xor_58_nl
      , loop_DES_rounds_5_xor_59_nl , loop_DES_rounds_5_xor_60_nl};
  wire[0:0] loop_DES_rounds_5_xor_44_nl;
  wire[0:0] loop_DES_rounds_5_xor_49_nl;
  wire[0:0] loop_DES_rounds_5_xor_45_nl;
  wire[0:0] loop_DES_rounds_5_xor_46_nl;
  wire[0:0] loop_DES_rounds_5_xor_47_nl;
  wire[0:0] loop_DES_rounds_5_xor_48_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_36_rg_addr;
  assign loop_DES_rounds_5_xor_44_nl = R_24_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_5_xor_49_nl = R_19_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_5_xor_45_nl = R_23_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_5_xor_46_nl = R_22_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign loop_DES_rounds_5_xor_47_nl = R_21_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_5_xor_48_nl = R_20_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_36_rg_addr = {3'b010 , loop_DES_rounds_5_xor_44_nl
      , loop_DES_rounds_5_xor_49_nl , loop_DES_rounds_5_xor_45_nl , loop_DES_rounds_5_xor_46_nl
      , loop_DES_rounds_5_xor_47_nl , loop_DES_rounds_5_xor_48_nl};
  wire[0:0] loop_DES_rounds_5_xor_62_nl;
  wire[0:0] loop_DES_rounds_5_xor_67_nl;
  wire[0:0] loop_DES_rounds_5_xor_63_nl;
  wire[0:0] loop_DES_rounds_5_xor_64_nl;
  wire[0:0] loop_DES_rounds_5_xor_65_nl;
  wire[0:0] loop_DES_rounds_5_xor_66_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_35_rg_addr;
  assign loop_DES_rounds_5_xor_62_nl = R_12_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_5_xor_67_nl = R_7_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_5_xor_63_nl = R_11_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_5_xor_64_nl = R_10_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_5_xor_65_nl = R_9_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_5_xor_66_nl = R_8_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_35_rg_addr = {3'b101 , loop_DES_rounds_5_xor_62_nl
      , loop_DES_rounds_5_xor_67_nl , loop_DES_rounds_5_xor_63_nl , loop_DES_rounds_5_xor_64_nl
      , loop_DES_rounds_5_xor_65_nl , loop_DES_rounds_5_xor_66_nl};
  wire[0:0] loop_DES_rounds_5_xor_74_nl;
  wire[0:0] loop_DES_rounds_5_xor_79_nl;
  wire[0:0] loop_DES_rounds_5_xor_75_nl;
  wire[0:0] loop_DES_rounds_5_xor_76_nl;
  wire[0:0] loop_DES_rounds_5_xor_77_nl;
  wire[0:0] loop_DES_rounds_5_xor_78_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_39_rg_addr;
  assign loop_DES_rounds_5_xor_74_nl = R_4_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_5_xor_79_nl = R_31_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign loop_DES_rounds_5_xor_75_nl = R_3_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_5_xor_76_nl = R_2_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_5_xor_77_nl = R_1_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_5_xor_78_nl = R_0_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_39_rg_addr = {3'b111 , loop_DES_rounds_5_xor_74_nl
      , loop_DES_rounds_5_xor_79_nl , loop_DES_rounds_5_xor_75_nl , loop_DES_rounds_5_xor_76_nl
      , loop_DES_rounds_5_xor_77_nl , loop_DES_rounds_5_xor_78_nl};
  wire[0:0] loop_DES_rounds_6_xor_50_nl;
  wire[0:0] loop_DES_rounds_6_xor_55_nl;
  wire[0:0] loop_DES_rounds_6_xor_51_nl;
  wire[0:0] loop_DES_rounds_6_xor_52_nl;
  wire[0:0] loop_DES_rounds_6_xor_53_nl;
  wire[0:0] loop_DES_rounds_6_xor_54_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_46_rg_addr;
  assign loop_DES_rounds_6_xor_50_nl = R_20_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_6_xor_55_nl = R_15_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_6_xor_51_nl = R_19_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign loop_DES_rounds_6_xor_52_nl = R_18_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_6_xor_53_nl = R_17_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign loop_DES_rounds_6_xor_54_nl = R_16_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_46_rg_addr = {3'b011 , loop_DES_rounds_6_xor_50_nl
      , loop_DES_rounds_6_xor_55_nl , loop_DES_rounds_6_xor_51_nl , loop_DES_rounds_6_xor_52_nl
      , loop_DES_rounds_6_xor_53_nl , loop_DES_rounds_6_xor_54_nl};
  wire[0:0] loop_DES_rounds_6_xor_68_nl;
  wire[0:0] loop_DES_rounds_6_xor_73_nl;
  wire[0:0] loop_DES_rounds_6_xor_69_nl;
  wire[0:0] loop_DES_rounds_6_xor_70_nl;
  wire[0:0] loop_DES_rounds_6_xor_71_nl;
  wire[0:0] loop_DES_rounds_6_xor_72_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_45_rg_addr;
  assign loop_DES_rounds_6_xor_68_nl = R_8_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_6_xor_73_nl = R_3_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_6_xor_69_nl = R_7_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_6_xor_70_nl = R_6_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_6_xor_71_nl = R_5_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_6_xor_72_nl = R_4_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_45_rg_addr = {3'b110 , loop_DES_rounds_6_xor_68_nl
      , loop_DES_rounds_6_xor_73_nl , loop_DES_rounds_6_xor_69_nl , loop_DES_rounds_6_xor_70_nl
      , loop_DES_rounds_6_xor_71_nl , loop_DES_rounds_6_xor_72_nl};
  wire[0:0] loop_DES_rounds_6_xor_38_nl;
  wire[0:0] loop_DES_rounds_6_xor_43_nl;
  wire[0:0] loop_DES_rounds_6_xor_39_nl;
  wire[0:0] loop_DES_rounds_6_xor_40_nl;
  wire[0:0] loop_DES_rounds_6_xor_41_nl;
  wire[0:0] loop_DES_rounds_6_xor_42_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_42_rg_addr;
  assign loop_DES_rounds_6_xor_38_nl = R_28_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign loop_DES_rounds_6_xor_43_nl = R_23_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign loop_DES_rounds_6_xor_39_nl = R_27_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_6_xor_40_nl = R_26_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_6_xor_41_nl = R_25_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_6_xor_42_nl = R_24_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_42_rg_addr = {3'b001 , loop_DES_rounds_6_xor_38_nl
      , loop_DES_rounds_6_xor_43_nl , loop_DES_rounds_6_xor_39_nl , loop_DES_rounds_6_xor_40_nl
      , loop_DES_rounds_6_xor_41_nl , loop_DES_rounds_6_xor_42_nl};
  wire[0:0] loop_DES_rounds_6_xor_nl;
  wire[0:0] loop_DES_rounds_6_xor_37_nl;
  wire[0:0] loop_DES_rounds_6_xor_33_nl;
  wire[0:0] loop_DES_rounds_6_xor_34_nl;
  wire[0:0] loop_DES_rounds_6_xor_35_nl;
  wire[0:0] loop_DES_rounds_6_xor_36_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_40_rg_addr;
  assign loop_DES_rounds_6_xor_nl = R_0_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_6_xor_37_nl = R_27_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign loop_DES_rounds_6_xor_33_nl = R_31_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_6_xor_34_nl = R_30_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_6_xor_35_nl = R_29_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_6_xor_36_nl = R_28_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_40_rg_addr = {3'b000 , loop_DES_rounds_6_xor_nl
      , loop_DES_rounds_6_xor_37_nl , loop_DES_rounds_6_xor_33_nl , loop_DES_rounds_6_xor_34_nl
      , loop_DES_rounds_6_xor_35_nl , loop_DES_rounds_6_xor_36_nl};
  wire[0:0] loop_DES_rounds_6_xor_56_nl;
  wire[0:0] loop_DES_rounds_6_xor_61_nl;
  wire[0:0] loop_DES_rounds_6_xor_57_nl;
  wire[0:0] loop_DES_rounds_6_xor_58_nl;
  wire[0:0] loop_DES_rounds_6_xor_59_nl;
  wire[0:0] loop_DES_rounds_6_xor_60_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_41_rg_addr;
  assign loop_DES_rounds_6_xor_56_nl = R_16_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_6_xor_61_nl = R_11_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_6_xor_57_nl = R_15_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_6_xor_58_nl = R_14_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_6_xor_59_nl = R_13_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_6_xor_60_nl = R_12_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_41_rg_addr = {3'b100 , loop_DES_rounds_6_xor_56_nl
      , loop_DES_rounds_6_xor_61_nl , loop_DES_rounds_6_xor_57_nl , loop_DES_rounds_6_xor_58_nl
      , loop_DES_rounds_6_xor_59_nl , loop_DES_rounds_6_xor_60_nl};
  wire[0:0] loop_DES_rounds_6_xor_44_nl;
  wire[0:0] loop_DES_rounds_6_xor_49_nl;
  wire[0:0] loop_DES_rounds_6_xor_45_nl;
  wire[0:0] loop_DES_rounds_6_xor_46_nl;
  wire[0:0] loop_DES_rounds_6_xor_47_nl;
  wire[0:0] loop_DES_rounds_6_xor_48_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_44_rg_addr;
  assign loop_DES_rounds_6_xor_44_nl = R_24_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_6_xor_49_nl = R_19_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_6_xor_45_nl = R_23_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_6_xor_46_nl = R_22_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_6_xor_47_nl = R_21_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_6_xor_48_nl = R_20_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_44_rg_addr = {3'b010 , loop_DES_rounds_6_xor_44_nl
      , loop_DES_rounds_6_xor_49_nl , loop_DES_rounds_6_xor_45_nl , loop_DES_rounds_6_xor_46_nl
      , loop_DES_rounds_6_xor_47_nl , loop_DES_rounds_6_xor_48_nl};
  wire[0:0] loop_DES_rounds_6_xor_62_nl;
  wire[0:0] loop_DES_rounds_6_xor_67_nl;
  wire[0:0] loop_DES_rounds_6_xor_63_nl;
  wire[0:0] loop_DES_rounds_6_xor_64_nl;
  wire[0:0] loop_DES_rounds_6_xor_65_nl;
  wire[0:0] loop_DES_rounds_6_xor_66_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_43_rg_addr;
  assign loop_DES_rounds_6_xor_62_nl = R_12_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign loop_DES_rounds_6_xor_67_nl = R_7_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_6_xor_63_nl = R_11_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_6_xor_64_nl = R_10_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_6_xor_65_nl = R_9_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_6_xor_66_nl = R_8_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_43_rg_addr = {3'b101 , loop_DES_rounds_6_xor_62_nl
      , loop_DES_rounds_6_xor_67_nl , loop_DES_rounds_6_xor_63_nl , loop_DES_rounds_6_xor_64_nl
      , loop_DES_rounds_6_xor_65_nl , loop_DES_rounds_6_xor_66_nl};
  wire[0:0] loop_DES_rounds_6_xor_74_nl;
  wire[0:0] loop_DES_rounds_6_xor_79_nl;
  wire[0:0] loop_DES_rounds_6_xor_75_nl;
  wire[0:0] loop_DES_rounds_6_xor_76_nl;
  wire[0:0] loop_DES_rounds_6_xor_77_nl;
  wire[0:0] loop_DES_rounds_6_xor_78_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_47_rg_addr;
  assign loop_DES_rounds_6_xor_74_nl = R_4_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_6_xor_79_nl = R_31_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_6_xor_75_nl = R_3_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_6_xor_76_nl = R_2_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_6_xor_77_nl = R_1_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_6_xor_78_nl = R_0_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_47_rg_addr = {3'b111 , loop_DES_rounds_6_xor_74_nl
      , loop_DES_rounds_6_xor_79_nl , loop_DES_rounds_6_xor_75_nl , loop_DES_rounds_6_xor_76_nl
      , loop_DES_rounds_6_xor_77_nl , loop_DES_rounds_6_xor_78_nl};
  wire[0:0] loop_DES_rounds_7_xor_50_nl;
  wire[0:0] loop_DES_rounds_7_xor_55_nl;
  wire[0:0] loop_DES_rounds_7_xor_51_nl;
  wire[0:0] loop_DES_rounds_7_xor_52_nl;
  wire[0:0] loop_DES_rounds_7_xor_53_nl;
  wire[0:0] loop_DES_rounds_7_xor_54_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_54_rg_addr;
  assign loop_DES_rounds_7_xor_50_nl = R_20_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign loop_DES_rounds_7_xor_55_nl = R_15_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_7_xor_51_nl = R_19_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_7_xor_52_nl = R_18_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign loop_DES_rounds_7_xor_53_nl = R_17_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign loop_DES_rounds_7_xor_54_nl = R_16_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_54_rg_addr = {3'b011 , loop_DES_rounds_7_xor_50_nl
      , loop_DES_rounds_7_xor_55_nl , loop_DES_rounds_7_xor_51_nl , loop_DES_rounds_7_xor_52_nl
      , loop_DES_rounds_7_xor_53_nl , loop_DES_rounds_7_xor_54_nl};
  wire[0:0] loop_DES_rounds_7_xor_68_nl;
  wire[0:0] loop_DES_rounds_7_xor_73_nl;
  wire[0:0] loop_DES_rounds_7_xor_69_nl;
  wire[0:0] loop_DES_rounds_7_xor_70_nl;
  wire[0:0] loop_DES_rounds_7_xor_71_nl;
  wire[0:0] loop_DES_rounds_7_xor_72_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_53_rg_addr;
  assign loop_DES_rounds_7_xor_68_nl = R_8_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_7_xor_73_nl = R_3_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_7_xor_69_nl = R_7_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_7_xor_70_nl = R_6_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_7_xor_71_nl = R_5_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign loop_DES_rounds_7_xor_72_nl = R_4_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_53_rg_addr = {3'b110 , loop_DES_rounds_7_xor_68_nl
      , loop_DES_rounds_7_xor_73_nl , loop_DES_rounds_7_xor_69_nl , loop_DES_rounds_7_xor_70_nl
      , loop_DES_rounds_7_xor_71_nl , loop_DES_rounds_7_xor_72_nl};
  wire[0:0] loop_DES_rounds_7_xor_38_nl;
  wire[0:0] loop_DES_rounds_7_xor_43_nl;
  wire[0:0] loop_DES_rounds_7_xor_39_nl;
  wire[0:0] loop_DES_rounds_7_xor_40_nl;
  wire[0:0] loop_DES_rounds_7_xor_41_nl;
  wire[0:0] loop_DES_rounds_7_xor_42_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_50_rg_addr;
  assign loop_DES_rounds_7_xor_38_nl = R_28_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign loop_DES_rounds_7_xor_43_nl = R_23_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_7_xor_39_nl = R_27_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_7_xor_40_nl = R_26_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_7_xor_41_nl = R_25_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_7_xor_42_nl = R_24_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_50_rg_addr = {3'b001 , loop_DES_rounds_7_xor_38_nl
      , loop_DES_rounds_7_xor_43_nl , loop_DES_rounds_7_xor_39_nl , loop_DES_rounds_7_xor_40_nl
      , loop_DES_rounds_7_xor_41_nl , loop_DES_rounds_7_xor_42_nl};
  wire[0:0] loop_DES_rounds_7_xor_nl;
  wire[0:0] loop_DES_rounds_7_xor_37_nl;
  wire[0:0] loop_DES_rounds_7_xor_33_nl;
  wire[0:0] loop_DES_rounds_7_xor_34_nl;
  wire[0:0] loop_DES_rounds_7_xor_35_nl;
  wire[0:0] loop_DES_rounds_7_xor_36_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_48_rg_addr;
  assign loop_DES_rounds_7_xor_nl = R_0_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_7_xor_37_nl = R_27_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign loop_DES_rounds_7_xor_33_nl = R_31_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_7_xor_34_nl = R_30_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_7_xor_35_nl = R_29_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_7_xor_36_nl = R_28_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_48_rg_addr = {3'b000 , loop_DES_rounds_7_xor_nl
      , loop_DES_rounds_7_xor_37_nl , loop_DES_rounds_7_xor_33_nl , loop_DES_rounds_7_xor_34_nl
      , loop_DES_rounds_7_xor_35_nl , loop_DES_rounds_7_xor_36_nl};
  wire[0:0] loop_DES_rounds_7_xor_56_nl;
  wire[0:0] loop_DES_rounds_7_xor_61_nl;
  wire[0:0] loop_DES_rounds_7_xor_57_nl;
  wire[0:0] loop_DES_rounds_7_xor_58_nl;
  wire[0:0] loop_DES_rounds_7_xor_59_nl;
  wire[0:0] loop_DES_rounds_7_xor_60_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_49_rg_addr;
  assign loop_DES_rounds_7_xor_56_nl = R_16_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_7_xor_61_nl = R_11_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_7_xor_57_nl = R_15_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign loop_DES_rounds_7_xor_58_nl = R_14_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_7_xor_59_nl = R_13_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_7_xor_60_nl = R_12_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_49_rg_addr = {3'b100 , loop_DES_rounds_7_xor_56_nl
      , loop_DES_rounds_7_xor_61_nl , loop_DES_rounds_7_xor_57_nl , loop_DES_rounds_7_xor_58_nl
      , loop_DES_rounds_7_xor_59_nl , loop_DES_rounds_7_xor_60_nl};
  wire[0:0] loop_DES_rounds_7_xor_44_nl;
  wire[0:0] loop_DES_rounds_7_xor_49_nl;
  wire[0:0] loop_DES_rounds_7_xor_45_nl;
  wire[0:0] loop_DES_rounds_7_xor_46_nl;
  wire[0:0] loop_DES_rounds_7_xor_47_nl;
  wire[0:0] loop_DES_rounds_7_xor_48_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_52_rg_addr;
  assign loop_DES_rounds_7_xor_44_nl = R_24_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_7_xor_49_nl = R_19_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign loop_DES_rounds_7_xor_45_nl = R_23_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_7_xor_46_nl = R_22_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_7_xor_47_nl = R_21_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_7_xor_48_nl = R_20_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_52_rg_addr = {3'b010 , loop_DES_rounds_7_xor_44_nl
      , loop_DES_rounds_7_xor_49_nl , loop_DES_rounds_7_xor_45_nl , loop_DES_rounds_7_xor_46_nl
      , loop_DES_rounds_7_xor_47_nl , loop_DES_rounds_7_xor_48_nl};
  wire[0:0] loop_DES_rounds_7_xor_62_nl;
  wire[0:0] loop_DES_rounds_7_xor_67_nl;
  wire[0:0] loop_DES_rounds_7_xor_63_nl;
  wire[0:0] loop_DES_rounds_7_xor_64_nl;
  wire[0:0] loop_DES_rounds_7_xor_65_nl;
  wire[0:0] loop_DES_rounds_7_xor_66_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_51_rg_addr;
  assign loop_DES_rounds_7_xor_62_nl = R_12_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_7_xor_67_nl = R_7_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_7_xor_63_nl = R_11_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_7_xor_64_nl = R_10_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_7_xor_65_nl = R_9_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_7_xor_66_nl = R_8_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_51_rg_addr = {3'b101 , loop_DES_rounds_7_xor_62_nl
      , loop_DES_rounds_7_xor_67_nl , loop_DES_rounds_7_xor_63_nl , loop_DES_rounds_7_xor_64_nl
      , loop_DES_rounds_7_xor_65_nl , loop_DES_rounds_7_xor_66_nl};
  wire[0:0] loop_DES_rounds_7_xor_74_nl;
  wire[0:0] loop_DES_rounds_7_xor_79_nl;
  wire[0:0] loop_DES_rounds_7_xor_75_nl;
  wire[0:0] loop_DES_rounds_7_xor_76_nl;
  wire[0:0] loop_DES_rounds_7_xor_77_nl;
  wire[0:0] loop_DES_rounds_7_xor_78_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_55_rg_addr;
  assign loop_DES_rounds_7_xor_74_nl = R_4_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_7_xor_79_nl = R_31_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_7_xor_75_nl = R_3_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_7_xor_76_nl = R_2_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_7_xor_77_nl = R_1_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_7_xor_78_nl = R_0_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_55_rg_addr = {3'b111 , loop_DES_rounds_7_xor_74_nl
      , loop_DES_rounds_7_xor_79_nl , loop_DES_rounds_7_xor_75_nl , loop_DES_rounds_7_xor_76_nl
      , loop_DES_rounds_7_xor_77_nl , loop_DES_rounds_7_xor_78_nl};
  wire[0:0] loop_DES_rounds_8_xor_50_nl;
  wire[0:0] loop_DES_rounds_8_xor_55_nl;
  wire[0:0] loop_DES_rounds_8_xor_51_nl;
  wire[0:0] loop_DES_rounds_8_xor_52_nl;
  wire[0:0] loop_DES_rounds_8_xor_53_nl;
  wire[0:0] loop_DES_rounds_8_xor_54_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_62_rg_addr;
  assign loop_DES_rounds_8_xor_50_nl = R_20_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign loop_DES_rounds_8_xor_55_nl = R_15_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_8_xor_51_nl = R_19_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_8_xor_52_nl = R_18_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign loop_DES_rounds_8_xor_53_nl = R_17_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_8_xor_54_nl = R_16_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_62_rg_addr = {3'b011 , loop_DES_rounds_8_xor_50_nl
      , loop_DES_rounds_8_xor_55_nl , loop_DES_rounds_8_xor_51_nl , loop_DES_rounds_8_xor_52_nl
      , loop_DES_rounds_8_xor_53_nl , loop_DES_rounds_8_xor_54_nl};
  wire[0:0] loop_DES_rounds_8_xor_68_nl;
  wire[0:0] loop_DES_rounds_8_xor_73_nl;
  wire[0:0] loop_DES_rounds_8_xor_69_nl;
  wire[0:0] loop_DES_rounds_8_xor_70_nl;
  wire[0:0] loop_DES_rounds_8_xor_71_nl;
  wire[0:0] loop_DES_rounds_8_xor_72_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_61_rg_addr;
  assign loop_DES_rounds_8_xor_68_nl = R_8_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_8_xor_73_nl = R_3_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_8_xor_69_nl = R_7_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_8_xor_70_nl = R_6_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_8_xor_71_nl = R_5_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_8_xor_72_nl = R_4_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_61_rg_addr = {3'b110 , loop_DES_rounds_8_xor_68_nl
      , loop_DES_rounds_8_xor_73_nl , loop_DES_rounds_8_xor_69_nl , loop_DES_rounds_8_xor_70_nl
      , loop_DES_rounds_8_xor_71_nl , loop_DES_rounds_8_xor_72_nl};
  wire[0:0] loop_DES_rounds_8_xor_38_nl;
  wire[0:0] loop_DES_rounds_8_xor_43_nl;
  wire[0:0] loop_DES_rounds_8_xor_39_nl;
  wire[0:0] loop_DES_rounds_8_xor_40_nl;
  wire[0:0] loop_DES_rounds_8_xor_41_nl;
  wire[0:0] loop_DES_rounds_8_xor_42_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_58_rg_addr;
  assign loop_DES_rounds_8_xor_38_nl = R_28_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign loop_DES_rounds_8_xor_43_nl = R_23_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_8_xor_39_nl = R_27_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_8_xor_40_nl = R_26_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_8_xor_41_nl = R_25_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign loop_DES_rounds_8_xor_42_nl = R_24_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_58_rg_addr = {3'b001 , loop_DES_rounds_8_xor_38_nl
      , loop_DES_rounds_8_xor_43_nl , loop_DES_rounds_8_xor_39_nl , loop_DES_rounds_8_xor_40_nl
      , loop_DES_rounds_8_xor_41_nl , loop_DES_rounds_8_xor_42_nl};
  wire[0:0] loop_DES_rounds_8_xor_nl;
  wire[0:0] loop_DES_rounds_8_xor_37_nl;
  wire[0:0] loop_DES_rounds_8_xor_33_nl;
  wire[0:0] loop_DES_rounds_8_xor_34_nl;
  wire[0:0] loop_DES_rounds_8_xor_35_nl;
  wire[0:0] loop_DES_rounds_8_xor_36_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_56_rg_addr;
  assign loop_DES_rounds_8_xor_nl = R_0_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign loop_DES_rounds_8_xor_37_nl = R_27_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_8_xor_33_nl = R_31_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_8_xor_34_nl = R_30_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_8_xor_35_nl = R_29_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_8_xor_36_nl = R_28_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_56_rg_addr = {3'b000 , loop_DES_rounds_8_xor_nl
      , loop_DES_rounds_8_xor_37_nl , loop_DES_rounds_8_xor_33_nl , loop_DES_rounds_8_xor_34_nl
      , loop_DES_rounds_8_xor_35_nl , loop_DES_rounds_8_xor_36_nl};
  wire[0:0] loop_DES_rounds_8_xor_56_nl;
  wire[0:0] loop_DES_rounds_8_xor_61_nl;
  wire[0:0] loop_DES_rounds_8_xor_57_nl;
  wire[0:0] loop_DES_rounds_8_xor_58_nl;
  wire[0:0] loop_DES_rounds_8_xor_59_nl;
  wire[0:0] loop_DES_rounds_8_xor_60_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_57_rg_addr;
  assign loop_DES_rounds_8_xor_56_nl = R_16_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_8_xor_61_nl = R_11_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_8_xor_57_nl = R_15_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_8_xor_58_nl = R_14_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_8_xor_59_nl = R_13_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_8_xor_60_nl = R_12_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_57_rg_addr = {3'b100 , loop_DES_rounds_8_xor_56_nl
      , loop_DES_rounds_8_xor_61_nl , loop_DES_rounds_8_xor_57_nl , loop_DES_rounds_8_xor_58_nl
      , loop_DES_rounds_8_xor_59_nl , loop_DES_rounds_8_xor_60_nl};
  wire[0:0] loop_DES_rounds_8_xor_44_nl;
  wire[0:0] loop_DES_rounds_8_xor_49_nl;
  wire[0:0] loop_DES_rounds_8_xor_45_nl;
  wire[0:0] loop_DES_rounds_8_xor_46_nl;
  wire[0:0] loop_DES_rounds_8_xor_47_nl;
  wire[0:0] loop_DES_rounds_8_xor_48_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_60_rg_addr;
  assign loop_DES_rounds_8_xor_44_nl = R_24_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_8_xor_49_nl = R_19_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_8_xor_45_nl = R_23_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_8_xor_46_nl = R_22_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_8_xor_47_nl = R_21_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_8_xor_48_nl = R_20_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_60_rg_addr = {3'b010 , loop_DES_rounds_8_xor_44_nl
      , loop_DES_rounds_8_xor_49_nl , loop_DES_rounds_8_xor_45_nl , loop_DES_rounds_8_xor_46_nl
      , loop_DES_rounds_8_xor_47_nl , loop_DES_rounds_8_xor_48_nl};
  wire[0:0] loop_DES_rounds_8_xor_62_nl;
  wire[0:0] loop_DES_rounds_8_xor_67_nl;
  wire[0:0] loop_DES_rounds_8_xor_63_nl;
  wire[0:0] loop_DES_rounds_8_xor_64_nl;
  wire[0:0] loop_DES_rounds_8_xor_65_nl;
  wire[0:0] loop_DES_rounds_8_xor_66_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_59_rg_addr;
  assign loop_DES_rounds_8_xor_62_nl = R_12_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_8_xor_67_nl = R_7_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_8_xor_63_nl = R_11_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_8_xor_64_nl = R_10_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_8_xor_65_nl = R_9_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_8_xor_66_nl = R_8_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_59_rg_addr = {3'b101 , loop_DES_rounds_8_xor_62_nl
      , loop_DES_rounds_8_xor_67_nl , loop_DES_rounds_8_xor_63_nl , loop_DES_rounds_8_xor_64_nl
      , loop_DES_rounds_8_xor_65_nl , loop_DES_rounds_8_xor_66_nl};
  wire[0:0] loop_DES_rounds_8_xor_74_nl;
  wire[0:0] loop_DES_rounds_8_xor_79_nl;
  wire[0:0] loop_DES_rounds_8_xor_75_nl;
  wire[0:0] loop_DES_rounds_8_xor_76_nl;
  wire[0:0] loop_DES_rounds_8_xor_77_nl;
  wire[0:0] loop_DES_rounds_8_xor_78_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_63_rg_addr;
  assign loop_DES_rounds_8_xor_74_nl = R_4_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_8_xor_79_nl = R_31_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_8_xor_75_nl = R_3_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_8_xor_76_nl = R_2_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign loop_DES_rounds_8_xor_77_nl = R_1_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_8_xor_78_nl = R_0_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_63_rg_addr = {3'b111 , loop_DES_rounds_8_xor_74_nl
      , loop_DES_rounds_8_xor_79_nl , loop_DES_rounds_8_xor_75_nl , loop_DES_rounds_8_xor_76_nl
      , loop_DES_rounds_8_xor_77_nl , loop_DES_rounds_8_xor_78_nl};
  wire[0:0] loop_DES_rounds_9_xor_50_nl;
  wire[0:0] loop_DES_rounds_9_xor_55_nl;
  wire[0:0] loop_DES_rounds_9_xor_51_nl;
  wire[0:0] loop_DES_rounds_9_xor_52_nl;
  wire[0:0] loop_DES_rounds_9_xor_53_nl;
  wire[0:0] loop_DES_rounds_9_xor_54_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_70_rg_addr;
  assign loop_DES_rounds_9_xor_50_nl = R_20_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_9_xor_55_nl = R_15_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign loop_DES_rounds_9_xor_51_nl = R_19_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_9_xor_52_nl = R_18_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_9_xor_53_nl = R_17_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_9_xor_54_nl = R_16_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_70_rg_addr = {3'b011 , loop_DES_rounds_9_xor_50_nl
      , loop_DES_rounds_9_xor_55_nl , loop_DES_rounds_9_xor_51_nl , loop_DES_rounds_9_xor_52_nl
      , loop_DES_rounds_9_xor_53_nl , loop_DES_rounds_9_xor_54_nl};
  wire[0:0] loop_DES_rounds_9_xor_68_nl;
  wire[0:0] loop_DES_rounds_9_xor_73_nl;
  wire[0:0] loop_DES_rounds_9_xor_69_nl;
  wire[0:0] loop_DES_rounds_9_xor_70_nl;
  wire[0:0] loop_DES_rounds_9_xor_71_nl;
  wire[0:0] loop_DES_rounds_9_xor_72_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_69_rg_addr;
  assign loop_DES_rounds_9_xor_68_nl = R_8_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_9_xor_73_nl = R_3_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign loop_DES_rounds_9_xor_69_nl = R_7_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign loop_DES_rounds_9_xor_70_nl = R_6_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_9_xor_71_nl = R_5_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_9_xor_72_nl = R_4_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_69_rg_addr = {3'b110 , loop_DES_rounds_9_xor_68_nl
      , loop_DES_rounds_9_xor_73_nl , loop_DES_rounds_9_xor_69_nl , loop_DES_rounds_9_xor_70_nl
      , loop_DES_rounds_9_xor_71_nl , loop_DES_rounds_9_xor_72_nl};
  wire[0:0] loop_DES_rounds_9_xor_38_nl;
  wire[0:0] loop_DES_rounds_9_xor_43_nl;
  wire[0:0] loop_DES_rounds_9_xor_39_nl;
  wire[0:0] loop_DES_rounds_9_xor_40_nl;
  wire[0:0] loop_DES_rounds_9_xor_41_nl;
  wire[0:0] loop_DES_rounds_9_xor_42_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_66_rg_addr;
  assign loop_DES_rounds_9_xor_38_nl = R_28_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_9_xor_43_nl = R_23_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_9_xor_39_nl = R_27_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign loop_DES_rounds_9_xor_40_nl = R_26_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign loop_DES_rounds_9_xor_41_nl = R_25_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_9_xor_42_nl = R_24_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_66_rg_addr = {3'b001 , loop_DES_rounds_9_xor_38_nl
      , loop_DES_rounds_9_xor_43_nl , loop_DES_rounds_9_xor_39_nl , loop_DES_rounds_9_xor_40_nl
      , loop_DES_rounds_9_xor_41_nl , loop_DES_rounds_9_xor_42_nl};
  wire[0:0] loop_DES_rounds_9_xor_nl;
  wire[0:0] loop_DES_rounds_9_xor_37_nl;
  wire[0:0] loop_DES_rounds_9_xor_33_nl;
  wire[0:0] loop_DES_rounds_9_xor_34_nl;
  wire[0:0] loop_DES_rounds_9_xor_35_nl;
  wire[0:0] loop_DES_rounds_9_xor_36_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_64_rg_addr;
  assign loop_DES_rounds_9_xor_nl = R_0_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_9_xor_37_nl = R_27_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign loop_DES_rounds_9_xor_33_nl = R_31_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign loop_DES_rounds_9_xor_34_nl = R_30_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_9_xor_35_nl = R_29_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign loop_DES_rounds_9_xor_36_nl = R_28_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_64_rg_addr = {3'b000 , loop_DES_rounds_9_xor_nl
      , loop_DES_rounds_9_xor_37_nl , loop_DES_rounds_9_xor_33_nl , loop_DES_rounds_9_xor_34_nl
      , loop_DES_rounds_9_xor_35_nl , loop_DES_rounds_9_xor_36_nl};
  wire[0:0] loop_DES_rounds_9_xor_56_nl;
  wire[0:0] loop_DES_rounds_9_xor_61_nl;
  wire[0:0] loop_DES_rounds_9_xor_57_nl;
  wire[0:0] loop_DES_rounds_9_xor_58_nl;
  wire[0:0] loop_DES_rounds_9_xor_59_nl;
  wire[0:0] loop_DES_rounds_9_xor_60_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_65_rg_addr;
  assign loop_DES_rounds_9_xor_56_nl = R_16_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_9_xor_61_nl = R_11_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_9_xor_57_nl = R_15_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_9_xor_58_nl = R_14_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_9_xor_59_nl = R_13_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_9_xor_60_nl = R_12_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_65_rg_addr = {3'b100 , loop_DES_rounds_9_xor_56_nl
      , loop_DES_rounds_9_xor_61_nl , loop_DES_rounds_9_xor_57_nl , loop_DES_rounds_9_xor_58_nl
      , loop_DES_rounds_9_xor_59_nl , loop_DES_rounds_9_xor_60_nl};
  wire[0:0] loop_DES_rounds_9_xor_44_nl;
  wire[0:0] loop_DES_rounds_9_xor_49_nl;
  wire[0:0] loop_DES_rounds_9_xor_45_nl;
  wire[0:0] loop_DES_rounds_9_xor_46_nl;
  wire[0:0] loop_DES_rounds_9_xor_47_nl;
  wire[0:0] loop_DES_rounds_9_xor_48_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_68_rg_addr;
  assign loop_DES_rounds_9_xor_44_nl = R_24_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_9_xor_49_nl = R_19_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_9_xor_45_nl = R_23_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_9_xor_46_nl = R_22_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_9_xor_47_nl = R_21_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_9_xor_48_nl = R_20_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_68_rg_addr = {3'b010 , loop_DES_rounds_9_xor_44_nl
      , loop_DES_rounds_9_xor_49_nl , loop_DES_rounds_9_xor_45_nl , loop_DES_rounds_9_xor_46_nl
      , loop_DES_rounds_9_xor_47_nl , loop_DES_rounds_9_xor_48_nl};
  wire[0:0] loop_DES_rounds_9_xor_62_nl;
  wire[0:0] loop_DES_rounds_9_xor_67_nl;
  wire[0:0] loop_DES_rounds_9_xor_63_nl;
  wire[0:0] loop_DES_rounds_9_xor_64_nl;
  wire[0:0] loop_DES_rounds_9_xor_65_nl;
  wire[0:0] loop_DES_rounds_9_xor_66_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_67_rg_addr;
  assign loop_DES_rounds_9_xor_62_nl = R_12_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_9_xor_67_nl = R_7_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_9_xor_63_nl = R_11_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_9_xor_64_nl = R_10_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_9_xor_65_nl = R_9_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_9_xor_66_nl = R_8_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_67_rg_addr = {3'b101 , loop_DES_rounds_9_xor_62_nl
      , loop_DES_rounds_9_xor_67_nl , loop_DES_rounds_9_xor_63_nl , loop_DES_rounds_9_xor_64_nl
      , loop_DES_rounds_9_xor_65_nl , loop_DES_rounds_9_xor_66_nl};
  wire[0:0] loop_DES_rounds_9_xor_74_nl;
  wire[0:0] loop_DES_rounds_9_xor_79_nl;
  wire[0:0] loop_DES_rounds_9_xor_75_nl;
  wire[0:0] loop_DES_rounds_9_xor_76_nl;
  wire[0:0] loop_DES_rounds_9_xor_77_nl;
  wire[0:0] loop_DES_rounds_9_xor_78_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_71_rg_addr;
  assign loop_DES_rounds_9_xor_74_nl = R_4_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_9_xor_79_nl = R_31_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_9_xor_75_nl = R_3_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_9_xor_76_nl = R_2_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_9_xor_77_nl = R_1_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_9_xor_78_nl = R_0_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_71_rg_addr = {3'b111 , loop_DES_rounds_9_xor_74_nl
      , loop_DES_rounds_9_xor_79_nl , loop_DES_rounds_9_xor_75_nl , loop_DES_rounds_9_xor_76_nl
      , loop_DES_rounds_9_xor_77_nl , loop_DES_rounds_9_xor_78_nl};
  wire[0:0] loop_DES_rounds_10_xor_50_nl;
  wire[0:0] loop_DES_rounds_10_xor_55_nl;
  wire[0:0] loop_DES_rounds_10_xor_51_nl;
  wire[0:0] loop_DES_rounds_10_xor_52_nl;
  wire[0:0] loop_DES_rounds_10_xor_53_nl;
  wire[0:0] loop_DES_rounds_10_xor_54_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_78_rg_addr;
  assign loop_DES_rounds_10_xor_50_nl = R_20_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_10_xor_55_nl = R_15_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_10_xor_51_nl = R_19_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_10_xor_52_nl = R_18_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_10_xor_53_nl = R_17_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_10_xor_54_nl = R_16_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_78_rg_addr = {3'b011 , loop_DES_rounds_10_xor_50_nl
      , loop_DES_rounds_10_xor_55_nl , loop_DES_rounds_10_xor_51_nl , loop_DES_rounds_10_xor_52_nl
      , loop_DES_rounds_10_xor_53_nl , loop_DES_rounds_10_xor_54_nl};
  wire[0:0] loop_DES_rounds_10_xor_68_nl;
  wire[0:0] loop_DES_rounds_10_xor_73_nl;
  wire[0:0] loop_DES_rounds_10_xor_69_nl;
  wire[0:0] loop_DES_rounds_10_xor_70_nl;
  wire[0:0] loop_DES_rounds_10_xor_71_nl;
  wire[0:0] loop_DES_rounds_10_xor_72_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_77_rg_addr;
  assign loop_DES_rounds_10_xor_68_nl = R_8_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_10_xor_73_nl = R_3_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_10_xor_69_nl = R_7_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_10_xor_70_nl = R_6_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_10_xor_71_nl = R_5_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_10_xor_72_nl = R_4_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_77_rg_addr = {3'b110 , loop_DES_rounds_10_xor_68_nl
      , loop_DES_rounds_10_xor_73_nl , loop_DES_rounds_10_xor_69_nl , loop_DES_rounds_10_xor_70_nl
      , loop_DES_rounds_10_xor_71_nl , loop_DES_rounds_10_xor_72_nl};
  wire[0:0] loop_DES_rounds_10_xor_38_nl;
  wire[0:0] loop_DES_rounds_10_xor_43_nl;
  wire[0:0] loop_DES_rounds_10_xor_39_nl;
  wire[0:0] loop_DES_rounds_10_xor_40_nl;
  wire[0:0] loop_DES_rounds_10_xor_41_nl;
  wire[0:0] loop_DES_rounds_10_xor_42_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_74_rg_addr;
  assign loop_DES_rounds_10_xor_38_nl = R_28_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign loop_DES_rounds_10_xor_43_nl = R_23_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_10_xor_39_nl = R_27_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign loop_DES_rounds_10_xor_40_nl = R_26_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign loop_DES_rounds_10_xor_41_nl = R_25_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_10_xor_42_nl = R_24_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_74_rg_addr = {3'b001 , loop_DES_rounds_10_xor_38_nl
      , loop_DES_rounds_10_xor_43_nl , loop_DES_rounds_10_xor_39_nl , loop_DES_rounds_10_xor_40_nl
      , loop_DES_rounds_10_xor_41_nl , loop_DES_rounds_10_xor_42_nl};
  wire[0:0] loop_DES_rounds_10_xor_nl;
  wire[0:0] loop_DES_rounds_10_xor_37_nl;
  wire[0:0] loop_DES_rounds_10_xor_33_nl;
  wire[0:0] loop_DES_rounds_10_xor_34_nl;
  wire[0:0] loop_DES_rounds_10_xor_35_nl;
  wire[0:0] loop_DES_rounds_10_xor_36_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_72_rg_addr;
  assign loop_DES_rounds_10_xor_nl = R_0_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_10_xor_37_nl = R_27_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_10_xor_33_nl = R_31_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_10_xor_34_nl = R_30_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign loop_DES_rounds_10_xor_35_nl = R_29_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign loop_DES_rounds_10_xor_36_nl = R_28_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_72_rg_addr = {3'b000 , loop_DES_rounds_10_xor_nl
      , loop_DES_rounds_10_xor_37_nl , loop_DES_rounds_10_xor_33_nl , loop_DES_rounds_10_xor_34_nl
      , loop_DES_rounds_10_xor_35_nl , loop_DES_rounds_10_xor_36_nl};
  wire[0:0] loop_DES_rounds_10_xor_56_nl;
  wire[0:0] loop_DES_rounds_10_xor_61_nl;
  wire[0:0] loop_DES_rounds_10_xor_57_nl;
  wire[0:0] loop_DES_rounds_10_xor_58_nl;
  wire[0:0] loop_DES_rounds_10_xor_59_nl;
  wire[0:0] loop_DES_rounds_10_xor_60_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_73_rg_addr;
  assign loop_DES_rounds_10_xor_56_nl = R_16_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_10_xor_61_nl = R_11_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_10_xor_57_nl = R_15_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_10_xor_58_nl = R_14_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_10_xor_59_nl = R_13_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_10_xor_60_nl = R_12_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_73_rg_addr = {3'b100 , loop_DES_rounds_10_xor_56_nl
      , loop_DES_rounds_10_xor_61_nl , loop_DES_rounds_10_xor_57_nl , loop_DES_rounds_10_xor_58_nl
      , loop_DES_rounds_10_xor_59_nl , loop_DES_rounds_10_xor_60_nl};
  wire[0:0] loop_DES_rounds_10_xor_44_nl;
  wire[0:0] loop_DES_rounds_10_xor_49_nl;
  wire[0:0] loop_DES_rounds_10_xor_45_nl;
  wire[0:0] loop_DES_rounds_10_xor_46_nl;
  wire[0:0] loop_DES_rounds_10_xor_47_nl;
  wire[0:0] loop_DES_rounds_10_xor_48_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_76_rg_addr;
  assign loop_DES_rounds_10_xor_44_nl = R_24_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_10_xor_49_nl = R_19_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_10_xor_45_nl = R_23_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_10_xor_46_nl = R_22_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_10_xor_47_nl = R_21_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_10_xor_48_nl = R_20_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_76_rg_addr = {3'b010 , loop_DES_rounds_10_xor_44_nl
      , loop_DES_rounds_10_xor_49_nl , loop_DES_rounds_10_xor_45_nl , loop_DES_rounds_10_xor_46_nl
      , loop_DES_rounds_10_xor_47_nl , loop_DES_rounds_10_xor_48_nl};
  wire[0:0] loop_DES_rounds_10_xor_62_nl;
  wire[0:0] loop_DES_rounds_10_xor_67_nl;
  wire[0:0] loop_DES_rounds_10_xor_63_nl;
  wire[0:0] loop_DES_rounds_10_xor_64_nl;
  wire[0:0] loop_DES_rounds_10_xor_65_nl;
  wire[0:0] loop_DES_rounds_10_xor_66_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_75_rg_addr;
  assign loop_DES_rounds_10_xor_62_nl = R_12_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_10_xor_67_nl = R_7_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_10_xor_63_nl = R_11_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_10_xor_64_nl = R_10_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign loop_DES_rounds_10_xor_65_nl = R_9_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_10_xor_66_nl = R_8_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_75_rg_addr = {3'b101 , loop_DES_rounds_10_xor_62_nl
      , loop_DES_rounds_10_xor_67_nl , loop_DES_rounds_10_xor_63_nl , loop_DES_rounds_10_xor_64_nl
      , loop_DES_rounds_10_xor_65_nl , loop_DES_rounds_10_xor_66_nl};
  wire[0:0] loop_DES_rounds_10_xor_74_nl;
  wire[0:0] loop_DES_rounds_10_xor_79_nl;
  wire[0:0] loop_DES_rounds_10_xor_75_nl;
  wire[0:0] loop_DES_rounds_10_xor_76_nl;
  wire[0:0] loop_DES_rounds_10_xor_77_nl;
  wire[0:0] loop_DES_rounds_10_xor_78_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_79_rg_addr;
  assign loop_DES_rounds_10_xor_74_nl = R_4_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_10_xor_79_nl = R_31_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_10_xor_75_nl = R_3_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_10_xor_76_nl = R_2_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_10_xor_77_nl = R_1_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_10_xor_78_nl = R_0_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_79_rg_addr = {3'b111 , loop_DES_rounds_10_xor_74_nl
      , loop_DES_rounds_10_xor_79_nl , loop_DES_rounds_10_xor_75_nl , loop_DES_rounds_10_xor_76_nl
      , loop_DES_rounds_10_xor_77_nl , loop_DES_rounds_10_xor_78_nl};
  wire[0:0] loop_DES_rounds_11_xor_50_nl;
  wire[0:0] loop_DES_rounds_11_xor_55_nl;
  wire[0:0] loop_DES_rounds_11_xor_51_nl;
  wire[0:0] loop_DES_rounds_11_xor_52_nl;
  wire[0:0] loop_DES_rounds_11_xor_53_nl;
  wire[0:0] loop_DES_rounds_11_xor_54_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_86_rg_addr;
  assign loop_DES_rounds_11_xor_50_nl = R_20_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_11_xor_55_nl = R_15_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_11_xor_51_nl = R_19_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_11_xor_52_nl = R_18_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_11_xor_53_nl = R_17_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign loop_DES_rounds_11_xor_54_nl = R_16_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_86_rg_addr = {3'b011 , loop_DES_rounds_11_xor_50_nl
      , loop_DES_rounds_11_xor_55_nl , loop_DES_rounds_11_xor_51_nl , loop_DES_rounds_11_xor_52_nl
      , loop_DES_rounds_11_xor_53_nl , loop_DES_rounds_11_xor_54_nl};
  wire[0:0] loop_DES_rounds_11_xor_68_nl;
  wire[0:0] loop_DES_rounds_11_xor_73_nl;
  wire[0:0] loop_DES_rounds_11_xor_69_nl;
  wire[0:0] loop_DES_rounds_11_xor_70_nl;
  wire[0:0] loop_DES_rounds_11_xor_71_nl;
  wire[0:0] loop_DES_rounds_11_xor_72_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_85_rg_addr;
  assign loop_DES_rounds_11_xor_68_nl = R_8_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_11_xor_73_nl = R_3_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_11_xor_69_nl = R_7_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign loop_DES_rounds_11_xor_70_nl = R_6_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_11_xor_71_nl = R_5_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_11_xor_72_nl = R_4_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_85_rg_addr = {3'b110 , loop_DES_rounds_11_xor_68_nl
      , loop_DES_rounds_11_xor_73_nl , loop_DES_rounds_11_xor_69_nl , loop_DES_rounds_11_xor_70_nl
      , loop_DES_rounds_11_xor_71_nl , loop_DES_rounds_11_xor_72_nl};
  wire[0:0] loop_DES_rounds_11_xor_38_nl;
  wire[0:0] loop_DES_rounds_11_xor_43_nl;
  wire[0:0] loop_DES_rounds_11_xor_39_nl;
  wire[0:0] loop_DES_rounds_11_xor_40_nl;
  wire[0:0] loop_DES_rounds_11_xor_41_nl;
  wire[0:0] loop_DES_rounds_11_xor_42_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_82_rg_addr;
  assign loop_DES_rounds_11_xor_38_nl = R_28_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_11_xor_43_nl = R_23_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_11_xor_39_nl = R_27_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_11_xor_40_nl = R_26_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_11_xor_41_nl = R_25_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_11_xor_42_nl = R_24_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_82_rg_addr = {3'b001 , loop_DES_rounds_11_xor_38_nl
      , loop_DES_rounds_11_xor_43_nl , loop_DES_rounds_11_xor_39_nl , loop_DES_rounds_11_xor_40_nl
      , loop_DES_rounds_11_xor_41_nl , loop_DES_rounds_11_xor_42_nl};
  wire[0:0] loop_DES_rounds_11_xor_nl;
  wire[0:0] loop_DES_rounds_11_xor_37_nl;
  wire[0:0] loop_DES_rounds_11_xor_33_nl;
  wire[0:0] loop_DES_rounds_11_xor_34_nl;
  wire[0:0] loop_DES_rounds_11_xor_35_nl;
  wire[0:0] loop_DES_rounds_11_xor_36_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_80_rg_addr;
  assign loop_DES_rounds_11_xor_nl = R_0_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_11_xor_37_nl = R_27_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_11_xor_33_nl = R_31_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_11_xor_34_nl = R_30_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign loop_DES_rounds_11_xor_35_nl = R_29_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign loop_DES_rounds_11_xor_36_nl = R_28_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_80_rg_addr = {3'b000 , loop_DES_rounds_11_xor_nl
      , loop_DES_rounds_11_xor_37_nl , loop_DES_rounds_11_xor_33_nl , loop_DES_rounds_11_xor_34_nl
      , loop_DES_rounds_11_xor_35_nl , loop_DES_rounds_11_xor_36_nl};
  wire[0:0] loop_DES_rounds_11_xor_56_nl;
  wire[0:0] loop_DES_rounds_11_xor_61_nl;
  wire[0:0] loop_DES_rounds_11_xor_57_nl;
  wire[0:0] loop_DES_rounds_11_xor_58_nl;
  wire[0:0] loop_DES_rounds_11_xor_59_nl;
  wire[0:0] loop_DES_rounds_11_xor_60_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_81_rg_addr;
  assign loop_DES_rounds_11_xor_56_nl = R_16_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_11_xor_61_nl = R_11_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_11_xor_57_nl = R_15_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_11_xor_58_nl = R_14_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_11_xor_59_nl = R_13_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_11_xor_60_nl = R_12_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_81_rg_addr = {3'b100 , loop_DES_rounds_11_xor_56_nl
      , loop_DES_rounds_11_xor_61_nl , loop_DES_rounds_11_xor_57_nl , loop_DES_rounds_11_xor_58_nl
      , loop_DES_rounds_11_xor_59_nl , loop_DES_rounds_11_xor_60_nl};
  wire[0:0] loop_DES_rounds_11_xor_44_nl;
  wire[0:0] loop_DES_rounds_11_xor_49_nl;
  wire[0:0] loop_DES_rounds_11_xor_45_nl;
  wire[0:0] loop_DES_rounds_11_xor_46_nl;
  wire[0:0] loop_DES_rounds_11_xor_47_nl;
  wire[0:0] loop_DES_rounds_11_xor_48_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_84_rg_addr;
  assign loop_DES_rounds_11_xor_44_nl = R_24_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_11_xor_49_nl = R_19_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_11_xor_45_nl = R_23_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_11_xor_46_nl = R_22_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_11_xor_47_nl = R_21_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_11_xor_48_nl = R_20_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_84_rg_addr = {3'b010 , loop_DES_rounds_11_xor_44_nl
      , loop_DES_rounds_11_xor_49_nl , loop_DES_rounds_11_xor_45_nl , loop_DES_rounds_11_xor_46_nl
      , loop_DES_rounds_11_xor_47_nl , loop_DES_rounds_11_xor_48_nl};
  wire[0:0] loop_DES_rounds_11_xor_62_nl;
  wire[0:0] loop_DES_rounds_11_xor_67_nl;
  wire[0:0] loop_DES_rounds_11_xor_63_nl;
  wire[0:0] loop_DES_rounds_11_xor_64_nl;
  wire[0:0] loop_DES_rounds_11_xor_65_nl;
  wire[0:0] loop_DES_rounds_11_xor_66_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_83_rg_addr;
  assign loop_DES_rounds_11_xor_62_nl = R_12_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_11_xor_67_nl = R_7_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_11_xor_63_nl = R_11_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_11_xor_64_nl = R_10_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_11_xor_65_nl = R_9_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign loop_DES_rounds_11_xor_66_nl = R_8_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_83_rg_addr = {3'b101 , loop_DES_rounds_11_xor_62_nl
      , loop_DES_rounds_11_xor_67_nl , loop_DES_rounds_11_xor_63_nl , loop_DES_rounds_11_xor_64_nl
      , loop_DES_rounds_11_xor_65_nl , loop_DES_rounds_11_xor_66_nl};
  wire[0:0] loop_DES_rounds_11_xor_74_nl;
  wire[0:0] loop_DES_rounds_11_xor_79_nl;
  wire[0:0] loop_DES_rounds_11_xor_75_nl;
  wire[0:0] loop_DES_rounds_11_xor_76_nl;
  wire[0:0] loop_DES_rounds_11_xor_77_nl;
  wire[0:0] loop_DES_rounds_11_xor_78_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_87_rg_addr;
  assign loop_DES_rounds_11_xor_74_nl = R_4_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_11_xor_79_nl = R_31_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_11_xor_75_nl = R_3_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_11_xor_76_nl = R_2_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_11_xor_77_nl = R_1_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_11_xor_78_nl = R_0_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_87_rg_addr = {3'b111 , loop_DES_rounds_11_xor_74_nl
      , loop_DES_rounds_11_xor_79_nl , loop_DES_rounds_11_xor_75_nl , loop_DES_rounds_11_xor_76_nl
      , loop_DES_rounds_11_xor_77_nl , loop_DES_rounds_11_xor_78_nl};
  wire[0:0] loop_DES_rounds_12_xor_50_nl;
  wire[0:0] loop_DES_rounds_12_xor_55_nl;
  wire[0:0] loop_DES_rounds_12_xor_51_nl;
  wire[0:0] loop_DES_rounds_12_xor_52_nl;
  wire[0:0] loop_DES_rounds_12_xor_53_nl;
  wire[0:0] loop_DES_rounds_12_xor_54_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_94_rg_addr;
  assign loop_DES_rounds_12_xor_50_nl = R_20_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_12_xor_55_nl = R_15_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_12_xor_51_nl = R_19_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign loop_DES_rounds_12_xor_52_nl = R_18_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign loop_DES_rounds_12_xor_53_nl = R_17_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign loop_DES_rounds_12_xor_54_nl = R_16_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_94_rg_addr = {3'b011 , loop_DES_rounds_12_xor_50_nl
      , loop_DES_rounds_12_xor_55_nl , loop_DES_rounds_12_xor_51_nl , loop_DES_rounds_12_xor_52_nl
      , loop_DES_rounds_12_xor_53_nl , loop_DES_rounds_12_xor_54_nl};
  wire[0:0] loop_DES_rounds_12_xor_68_nl;
  wire[0:0] loop_DES_rounds_12_xor_73_nl;
  wire[0:0] loop_DES_rounds_12_xor_69_nl;
  wire[0:0] loop_DES_rounds_12_xor_70_nl;
  wire[0:0] loop_DES_rounds_12_xor_71_nl;
  wire[0:0] loop_DES_rounds_12_xor_72_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_93_rg_addr;
  assign loop_DES_rounds_12_xor_68_nl = R_8_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_12_xor_73_nl = R_3_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_12_xor_69_nl = R_7_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_12_xor_70_nl = R_6_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_12_xor_71_nl = R_5_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_12_xor_72_nl = R_4_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_93_rg_addr = {3'b110 , loop_DES_rounds_12_xor_68_nl
      , loop_DES_rounds_12_xor_73_nl , loop_DES_rounds_12_xor_69_nl , loop_DES_rounds_12_xor_70_nl
      , loop_DES_rounds_12_xor_71_nl , loop_DES_rounds_12_xor_72_nl};
  wire[0:0] loop_DES_rounds_12_xor_38_nl;
  wire[0:0] loop_DES_rounds_12_xor_43_nl;
  wire[0:0] loop_DES_rounds_12_xor_39_nl;
  wire[0:0] loop_DES_rounds_12_xor_40_nl;
  wire[0:0] loop_DES_rounds_12_xor_41_nl;
  wire[0:0] loop_DES_rounds_12_xor_42_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_90_rg_addr;
  assign loop_DES_rounds_12_xor_38_nl = R_28_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_12_xor_43_nl = R_23_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_12_xor_39_nl = R_27_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_12_xor_40_nl = R_26_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_12_xor_41_nl = R_25_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_12_xor_42_nl = R_24_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_90_rg_addr = {3'b001 , loop_DES_rounds_12_xor_38_nl
      , loop_DES_rounds_12_xor_43_nl , loop_DES_rounds_12_xor_39_nl , loop_DES_rounds_12_xor_40_nl
      , loop_DES_rounds_12_xor_41_nl , loop_DES_rounds_12_xor_42_nl};
  wire[0:0] loop_DES_rounds_12_xor_nl;
  wire[0:0] loop_DES_rounds_12_xor_37_nl;
  wire[0:0] loop_DES_rounds_12_xor_33_nl;
  wire[0:0] loop_DES_rounds_12_xor_34_nl;
  wire[0:0] loop_DES_rounds_12_xor_35_nl;
  wire[0:0] loop_DES_rounds_12_xor_36_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_88_rg_addr;
  assign loop_DES_rounds_12_xor_nl = R_0_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_12_xor_37_nl = R_27_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_12_xor_33_nl = R_31_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_12_xor_34_nl = R_30_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign loop_DES_rounds_12_xor_35_nl = R_29_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign loop_DES_rounds_12_xor_36_nl = R_28_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_88_rg_addr = {3'b000 , loop_DES_rounds_12_xor_nl
      , loop_DES_rounds_12_xor_37_nl , loop_DES_rounds_12_xor_33_nl , loop_DES_rounds_12_xor_34_nl
      , loop_DES_rounds_12_xor_35_nl , loop_DES_rounds_12_xor_36_nl};
  wire[0:0] loop_DES_rounds_12_xor_56_nl;
  wire[0:0] loop_DES_rounds_12_xor_61_nl;
  wire[0:0] loop_DES_rounds_12_xor_57_nl;
  wire[0:0] loop_DES_rounds_12_xor_58_nl;
  wire[0:0] loop_DES_rounds_12_xor_59_nl;
  wire[0:0] loop_DES_rounds_12_xor_60_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_89_rg_addr;
  assign loop_DES_rounds_12_xor_56_nl = R_16_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_12_xor_61_nl = R_11_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_12_xor_57_nl = R_15_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_12_xor_58_nl = R_14_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_12_xor_59_nl = R_13_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_12_xor_60_nl = R_12_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_89_rg_addr = {3'b100 , loop_DES_rounds_12_xor_56_nl
      , loop_DES_rounds_12_xor_61_nl , loop_DES_rounds_12_xor_57_nl , loop_DES_rounds_12_xor_58_nl
      , loop_DES_rounds_12_xor_59_nl , loop_DES_rounds_12_xor_60_nl};
  wire[0:0] loop_DES_rounds_12_xor_44_nl;
  wire[0:0] loop_DES_rounds_12_xor_49_nl;
  wire[0:0] loop_DES_rounds_12_xor_45_nl;
  wire[0:0] loop_DES_rounds_12_xor_46_nl;
  wire[0:0] loop_DES_rounds_12_xor_47_nl;
  wire[0:0] loop_DES_rounds_12_xor_48_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_92_rg_addr;
  assign loop_DES_rounds_12_xor_44_nl = R_24_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_12_xor_49_nl = R_19_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_12_xor_45_nl = R_23_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_12_xor_46_nl = R_22_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_12_xor_47_nl = R_21_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_12_xor_48_nl = R_20_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_92_rg_addr = {3'b010 , loop_DES_rounds_12_xor_44_nl
      , loop_DES_rounds_12_xor_49_nl , loop_DES_rounds_12_xor_45_nl , loop_DES_rounds_12_xor_46_nl
      , loop_DES_rounds_12_xor_47_nl , loop_DES_rounds_12_xor_48_nl};
  wire[0:0] loop_DES_rounds_12_xor_62_nl;
  wire[0:0] loop_DES_rounds_12_xor_67_nl;
  wire[0:0] loop_DES_rounds_12_xor_63_nl;
  wire[0:0] loop_DES_rounds_12_xor_64_nl;
  wire[0:0] loop_DES_rounds_12_xor_65_nl;
  wire[0:0] loop_DES_rounds_12_xor_66_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_91_rg_addr;
  assign loop_DES_rounds_12_xor_62_nl = R_12_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_12_xor_67_nl = R_7_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_12_xor_63_nl = R_11_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_12_xor_64_nl = R_10_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_12_xor_65_nl = R_9_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_12_xor_66_nl = R_8_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_91_rg_addr = {3'b101 , loop_DES_rounds_12_xor_62_nl
      , loop_DES_rounds_12_xor_67_nl , loop_DES_rounds_12_xor_63_nl , loop_DES_rounds_12_xor_64_nl
      , loop_DES_rounds_12_xor_65_nl , loop_DES_rounds_12_xor_66_nl};
  wire[0:0] loop_DES_rounds_12_xor_74_nl;
  wire[0:0] loop_DES_rounds_12_xor_79_nl;
  wire[0:0] loop_DES_rounds_12_xor_75_nl;
  wire[0:0] loop_DES_rounds_12_xor_76_nl;
  wire[0:0] loop_DES_rounds_12_xor_77_nl;
  wire[0:0] loop_DES_rounds_12_xor_78_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_95_rg_addr;
  assign loop_DES_rounds_12_xor_74_nl = R_4_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_12_xor_79_nl = R_31_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_12_xor_75_nl = R_3_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_12_xor_76_nl = R_2_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_12_xor_77_nl = R_1_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_12_xor_78_nl = R_0_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_95_rg_addr = {3'b111 , loop_DES_rounds_12_xor_74_nl
      , loop_DES_rounds_12_xor_79_nl , loop_DES_rounds_12_xor_75_nl , loop_DES_rounds_12_xor_76_nl
      , loop_DES_rounds_12_xor_77_nl , loop_DES_rounds_12_xor_78_nl};
  wire[0:0] loop_DES_rounds_13_xor_50_nl;
  wire[0:0] loop_DES_rounds_13_xor_55_nl;
  wire[0:0] loop_DES_rounds_13_xor_51_nl;
  wire[0:0] loop_DES_rounds_13_xor_52_nl;
  wire[0:0] loop_DES_rounds_13_xor_53_nl;
  wire[0:0] loop_DES_rounds_13_xor_54_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_102_rg_addr;
  assign loop_DES_rounds_13_xor_50_nl = R_20_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign loop_DES_rounds_13_xor_55_nl = R_15_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_13_xor_51_nl = R_19_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign loop_DES_rounds_13_xor_52_nl = R_18_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_13_xor_53_nl = R_17_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign loop_DES_rounds_13_xor_54_nl = R_16_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_102_rg_addr = {3'b011 , loop_DES_rounds_13_xor_50_nl
      , loop_DES_rounds_13_xor_55_nl , loop_DES_rounds_13_xor_51_nl , loop_DES_rounds_13_xor_52_nl
      , loop_DES_rounds_13_xor_53_nl , loop_DES_rounds_13_xor_54_nl};
  wire[0:0] loop_DES_rounds_13_xor_68_nl;
  wire[0:0] loop_DES_rounds_13_xor_73_nl;
  wire[0:0] loop_DES_rounds_13_xor_69_nl;
  wire[0:0] loop_DES_rounds_13_xor_70_nl;
  wire[0:0] loop_DES_rounds_13_xor_71_nl;
  wire[0:0] loop_DES_rounds_13_xor_72_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_101_rg_addr;
  assign loop_DES_rounds_13_xor_68_nl = R_8_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_13_xor_73_nl = R_3_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_13_xor_69_nl = R_7_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_13_xor_70_nl = R_6_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_13_xor_71_nl = R_5_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_13_xor_72_nl = R_4_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_101_rg_addr = {3'b110 , loop_DES_rounds_13_xor_68_nl
      , loop_DES_rounds_13_xor_73_nl , loop_DES_rounds_13_xor_69_nl , loop_DES_rounds_13_xor_70_nl
      , loop_DES_rounds_13_xor_71_nl , loop_DES_rounds_13_xor_72_nl};
  wire[0:0] loop_DES_rounds_13_xor_38_nl;
  wire[0:0] loop_DES_rounds_13_xor_43_nl;
  wire[0:0] loop_DES_rounds_13_xor_39_nl;
  wire[0:0] loop_DES_rounds_13_xor_40_nl;
  wire[0:0] loop_DES_rounds_13_xor_41_nl;
  wire[0:0] loop_DES_rounds_13_xor_42_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_98_rg_addr;
  assign loop_DES_rounds_13_xor_38_nl = R_28_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_13_xor_43_nl = R_23_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_13_xor_39_nl = R_27_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_13_xor_40_nl = R_26_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_13_xor_41_nl = R_25_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_13_xor_42_nl = R_24_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_98_rg_addr = {3'b001 , loop_DES_rounds_13_xor_38_nl
      , loop_DES_rounds_13_xor_43_nl , loop_DES_rounds_13_xor_39_nl , loop_DES_rounds_13_xor_40_nl
      , loop_DES_rounds_13_xor_41_nl , loop_DES_rounds_13_xor_42_nl};
  wire[0:0] loop_DES_rounds_13_xor_nl;
  wire[0:0] loop_DES_rounds_13_xor_37_nl;
  wire[0:0] loop_DES_rounds_13_xor_33_nl;
  wire[0:0] loop_DES_rounds_13_xor_34_nl;
  wire[0:0] loop_DES_rounds_13_xor_35_nl;
  wire[0:0] loop_DES_rounds_13_xor_36_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_96_rg_addr;
  assign loop_DES_rounds_13_xor_nl = R_0_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_13_xor_37_nl = R_27_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign loop_DES_rounds_13_xor_33_nl = R_31_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_13_xor_34_nl = R_30_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_13_xor_35_nl = R_29_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_13_xor_36_nl = R_28_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_96_rg_addr = {3'b000 , loop_DES_rounds_13_xor_nl
      , loop_DES_rounds_13_xor_37_nl , loop_DES_rounds_13_xor_33_nl , loop_DES_rounds_13_xor_34_nl
      , loop_DES_rounds_13_xor_35_nl , loop_DES_rounds_13_xor_36_nl};
  wire[0:0] loop_DES_rounds_13_xor_56_nl;
  wire[0:0] loop_DES_rounds_13_xor_61_nl;
  wire[0:0] loop_DES_rounds_13_xor_57_nl;
  wire[0:0] loop_DES_rounds_13_xor_58_nl;
  wire[0:0] loop_DES_rounds_13_xor_59_nl;
  wire[0:0] loop_DES_rounds_13_xor_60_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_97_rg_addr;
  assign loop_DES_rounds_13_xor_56_nl = R_16_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign loop_DES_rounds_13_xor_61_nl = R_11_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_13_xor_57_nl = R_15_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_13_xor_58_nl = R_14_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_13_xor_59_nl = R_13_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_13_xor_60_nl = R_12_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_97_rg_addr = {3'b100 , loop_DES_rounds_13_xor_56_nl
      , loop_DES_rounds_13_xor_61_nl , loop_DES_rounds_13_xor_57_nl , loop_DES_rounds_13_xor_58_nl
      , loop_DES_rounds_13_xor_59_nl , loop_DES_rounds_13_xor_60_nl};
  wire[0:0] loop_DES_rounds_13_xor_44_nl;
  wire[0:0] loop_DES_rounds_13_xor_49_nl;
  wire[0:0] loop_DES_rounds_13_xor_45_nl;
  wire[0:0] loop_DES_rounds_13_xor_46_nl;
  wire[0:0] loop_DES_rounds_13_xor_47_nl;
  wire[0:0] loop_DES_rounds_13_xor_48_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_100_rg_addr;
  assign loop_DES_rounds_13_xor_44_nl = R_24_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_13_xor_49_nl = R_19_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_13_xor_45_nl = R_23_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_13_xor_46_nl = R_22_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_13_xor_47_nl = R_21_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_13_xor_48_nl = R_20_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_100_rg_addr = {3'b010 , loop_DES_rounds_13_xor_44_nl
      , loop_DES_rounds_13_xor_49_nl , loop_DES_rounds_13_xor_45_nl , loop_DES_rounds_13_xor_46_nl
      , loop_DES_rounds_13_xor_47_nl , loop_DES_rounds_13_xor_48_nl};
  wire[0:0] loop_DES_rounds_13_xor_62_nl;
  wire[0:0] loop_DES_rounds_13_xor_67_nl;
  wire[0:0] loop_DES_rounds_13_xor_63_nl;
  wire[0:0] loop_DES_rounds_13_xor_64_nl;
  wire[0:0] loop_DES_rounds_13_xor_65_nl;
  wire[0:0] loop_DES_rounds_13_xor_66_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_99_rg_addr;
  assign loop_DES_rounds_13_xor_62_nl = R_12_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_13_xor_67_nl = R_7_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_13_xor_63_nl = R_11_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_13_xor_64_nl = R_10_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_13_xor_65_nl = R_9_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign loop_DES_rounds_13_xor_66_nl = R_8_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_99_rg_addr = {3'b101 , loop_DES_rounds_13_xor_62_nl
      , loop_DES_rounds_13_xor_67_nl , loop_DES_rounds_13_xor_63_nl , loop_DES_rounds_13_xor_64_nl
      , loop_DES_rounds_13_xor_65_nl , loop_DES_rounds_13_xor_66_nl};
  wire[0:0] loop_DES_rounds_13_xor_74_nl;
  wire[0:0] loop_DES_rounds_13_xor_79_nl;
  wire[0:0] loop_DES_rounds_13_xor_75_nl;
  wire[0:0] loop_DES_rounds_13_xor_76_nl;
  wire[0:0] loop_DES_rounds_13_xor_77_nl;
  wire[0:0] loop_DES_rounds_13_xor_78_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_103_rg_addr;
  assign loop_DES_rounds_13_xor_74_nl = R_4_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_13_xor_79_nl = R_31_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_13_xor_75_nl = R_3_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_13_xor_76_nl = R_2_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_13_xor_77_nl = R_1_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_13_xor_78_nl = R_0_12_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_103_rg_addr = {3'b111 , loop_DES_rounds_13_xor_74_nl
      , loop_DES_rounds_13_xor_79_nl , loop_DES_rounds_13_xor_75_nl , loop_DES_rounds_13_xor_76_nl
      , loop_DES_rounds_13_xor_77_nl , loop_DES_rounds_13_xor_78_nl};
  wire[0:0] loop_DES_rounds_14_xor_50_nl;
  wire[0:0] loop_DES_rounds_14_xor_55_nl;
  wire[0:0] loop_DES_rounds_14_xor_51_nl;
  wire[0:0] loop_DES_rounds_14_xor_52_nl;
  wire[0:0] loop_DES_rounds_14_xor_53_nl;
  wire[0:0] loop_DES_rounds_14_xor_54_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_110_rg_addr;
  assign loop_DES_rounds_14_xor_50_nl = R_20_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign loop_DES_rounds_14_xor_55_nl = R_15_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_14_xor_51_nl = R_19_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign loop_DES_rounds_14_xor_52_nl = R_18_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_14_xor_53_nl = R_17_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign loop_DES_rounds_14_xor_54_nl = R_16_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_110_rg_addr = {3'b011 , loop_DES_rounds_14_xor_50_nl
      , loop_DES_rounds_14_xor_55_nl , loop_DES_rounds_14_xor_51_nl , loop_DES_rounds_14_xor_52_nl
      , loop_DES_rounds_14_xor_53_nl , loop_DES_rounds_14_xor_54_nl};
  wire[0:0] loop_DES_rounds_14_xor_68_nl;
  wire[0:0] loop_DES_rounds_14_xor_73_nl;
  wire[0:0] loop_DES_rounds_14_xor_69_nl;
  wire[0:0] loop_DES_rounds_14_xor_70_nl;
  wire[0:0] loop_DES_rounds_14_xor_71_nl;
  wire[0:0] loop_DES_rounds_14_xor_72_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_109_rg_addr;
  assign loop_DES_rounds_14_xor_68_nl = R_8_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_14_xor_73_nl = R_3_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_14_xor_69_nl = R_7_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_14_xor_70_nl = R_6_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign loop_DES_rounds_14_xor_71_nl = R_5_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_14_xor_72_nl = R_4_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_109_rg_addr = {3'b110 , loop_DES_rounds_14_xor_68_nl
      , loop_DES_rounds_14_xor_73_nl , loop_DES_rounds_14_xor_69_nl , loop_DES_rounds_14_xor_70_nl
      , loop_DES_rounds_14_xor_71_nl , loop_DES_rounds_14_xor_72_nl};
  wire[0:0] loop_DES_rounds_14_xor_38_nl;
  wire[0:0] loop_DES_rounds_14_xor_43_nl;
  wire[0:0] loop_DES_rounds_14_xor_39_nl;
  wire[0:0] loop_DES_rounds_14_xor_40_nl;
  wire[0:0] loop_DES_rounds_14_xor_41_nl;
  wire[0:0] loop_DES_rounds_14_xor_42_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_106_rg_addr;
  assign loop_DES_rounds_14_xor_38_nl = R_28_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign loop_DES_rounds_14_xor_43_nl = R_23_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_14_xor_39_nl = R_27_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_14_xor_40_nl = R_26_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_14_xor_41_nl = R_25_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_14_xor_42_nl = R_24_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_106_rg_addr = {3'b001 , loop_DES_rounds_14_xor_38_nl
      , loop_DES_rounds_14_xor_43_nl , loop_DES_rounds_14_xor_39_nl , loop_DES_rounds_14_xor_40_nl
      , loop_DES_rounds_14_xor_41_nl , loop_DES_rounds_14_xor_42_nl};
  wire[0:0] loop_DES_rounds_14_xor_nl;
  wire[0:0] loop_DES_rounds_14_xor_37_nl;
  wire[0:0] loop_DES_rounds_14_xor_33_nl;
  wire[0:0] loop_DES_rounds_14_xor_34_nl;
  wire[0:0] loop_DES_rounds_14_xor_35_nl;
  wire[0:0] loop_DES_rounds_14_xor_36_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_104_rg_addr;
  assign loop_DES_rounds_14_xor_nl = R_0_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign loop_DES_rounds_14_xor_37_nl = R_27_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign loop_DES_rounds_14_xor_33_nl = R_31_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_14_xor_34_nl = R_30_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_14_xor_35_nl = R_29_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_14_xor_36_nl = R_28_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_104_rg_addr = {3'b000 , loop_DES_rounds_14_xor_nl
      , loop_DES_rounds_14_xor_37_nl , loop_DES_rounds_14_xor_33_nl , loop_DES_rounds_14_xor_34_nl
      , loop_DES_rounds_14_xor_35_nl , loop_DES_rounds_14_xor_36_nl};
  wire[0:0] loop_DES_rounds_14_xor_56_nl;
  wire[0:0] loop_DES_rounds_14_xor_61_nl;
  wire[0:0] loop_DES_rounds_14_xor_57_nl;
  wire[0:0] loop_DES_rounds_14_xor_58_nl;
  wire[0:0] loop_DES_rounds_14_xor_59_nl;
  wire[0:0] loop_DES_rounds_14_xor_60_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_105_rg_addr;
  assign loop_DES_rounds_14_xor_56_nl = R_16_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_14_xor_61_nl = R_11_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_14_xor_57_nl = R_15_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_14_xor_58_nl = R_14_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_14_xor_59_nl = R_13_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_14_xor_60_nl = R_12_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_105_rg_addr = {3'b100 , loop_DES_rounds_14_xor_56_nl
      , loop_DES_rounds_14_xor_61_nl , loop_DES_rounds_14_xor_57_nl , loop_DES_rounds_14_xor_58_nl
      , loop_DES_rounds_14_xor_59_nl , loop_DES_rounds_14_xor_60_nl};
  wire[0:0] loop_DES_rounds_14_xor_44_nl;
  wire[0:0] loop_DES_rounds_14_xor_49_nl;
  wire[0:0] loop_DES_rounds_14_xor_45_nl;
  wire[0:0] loop_DES_rounds_14_xor_46_nl;
  wire[0:0] loop_DES_rounds_14_xor_47_nl;
  wire[0:0] loop_DES_rounds_14_xor_48_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_108_rg_addr;
  assign loop_DES_rounds_14_xor_44_nl = R_24_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign loop_DES_rounds_14_xor_49_nl = R_19_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_14_xor_45_nl = R_23_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_14_xor_46_nl = R_22_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_14_xor_47_nl = R_21_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_14_xor_48_nl = R_20_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_108_rg_addr = {3'b010 , loop_DES_rounds_14_xor_44_nl
      , loop_DES_rounds_14_xor_49_nl , loop_DES_rounds_14_xor_45_nl , loop_DES_rounds_14_xor_46_nl
      , loop_DES_rounds_14_xor_47_nl , loop_DES_rounds_14_xor_48_nl};
  wire[0:0] loop_DES_rounds_14_xor_62_nl;
  wire[0:0] loop_DES_rounds_14_xor_67_nl;
  wire[0:0] loop_DES_rounds_14_xor_63_nl;
  wire[0:0] loop_DES_rounds_14_xor_64_nl;
  wire[0:0] loop_DES_rounds_14_xor_65_nl;
  wire[0:0] loop_DES_rounds_14_xor_66_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_107_rg_addr;
  assign loop_DES_rounds_14_xor_62_nl = R_12_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_14_xor_67_nl = R_7_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_14_xor_63_nl = R_11_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_14_xor_64_nl = R_10_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_14_xor_65_nl = R_9_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_14_xor_66_nl = R_8_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_107_rg_addr = {3'b101 , loop_DES_rounds_14_xor_62_nl
      , loop_DES_rounds_14_xor_67_nl , loop_DES_rounds_14_xor_63_nl , loop_DES_rounds_14_xor_64_nl
      , loop_DES_rounds_14_xor_65_nl , loop_DES_rounds_14_xor_66_nl};
  wire[0:0] loop_DES_rounds_14_xor_74_nl;
  wire[0:0] loop_DES_rounds_14_xor_79_nl;
  wire[0:0] loop_DES_rounds_14_xor_75_nl;
  wire[0:0] loop_DES_rounds_14_xor_76_nl;
  wire[0:0] loop_DES_rounds_14_xor_77_nl;
  wire[0:0] loop_DES_rounds_14_xor_78_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_111_rg_addr;
  assign loop_DES_rounds_14_xor_74_nl = R_4_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_14_xor_79_nl = R_31_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_14_xor_75_nl = R_3_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_14_xor_76_nl = R_2_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_14_xor_77_nl = R_1_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_14_xor_78_nl = R_0_13_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_111_rg_addr = {3'b111 , loop_DES_rounds_14_xor_74_nl
      , loop_DES_rounds_14_xor_79_nl , loop_DES_rounds_14_xor_75_nl , loop_DES_rounds_14_xor_76_nl
      , loop_DES_rounds_14_xor_77_nl , loop_DES_rounds_14_xor_78_nl};
  wire[0:0] loop_DES_rounds_15_xor_50_nl;
  wire[0:0] loop_DES_rounds_15_xor_55_nl;
  wire[0:0] loop_DES_rounds_15_xor_51_nl;
  wire[0:0] loop_DES_rounds_15_xor_52_nl;
  wire[0:0] loop_DES_rounds_15_xor_53_nl;
  wire[0:0] loop_DES_rounds_15_xor_54_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_118_rg_addr;
  assign loop_DES_rounds_15_xor_50_nl = R_20_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign loop_DES_rounds_15_xor_55_nl = R_15_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_15_xor_51_nl = R_19_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_15_xor_52_nl = R_18_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_15_xor_53_nl = R_17_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_15_xor_54_nl = R_16_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_118_rg_addr = {3'b011 , loop_DES_rounds_15_xor_50_nl
      , loop_DES_rounds_15_xor_55_nl , loop_DES_rounds_15_xor_51_nl , loop_DES_rounds_15_xor_52_nl
      , loop_DES_rounds_15_xor_53_nl , loop_DES_rounds_15_xor_54_nl};
  wire[0:0] loop_DES_rounds_15_xor_68_nl;
  wire[0:0] loop_DES_rounds_15_xor_73_nl;
  wire[0:0] loop_DES_rounds_15_xor_69_nl;
  wire[0:0] loop_DES_rounds_15_xor_70_nl;
  wire[0:0] loop_DES_rounds_15_xor_71_nl;
  wire[0:0] loop_DES_rounds_15_xor_72_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_117_rg_addr;
  assign loop_DES_rounds_15_xor_68_nl = R_8_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_15_xor_73_nl = R_3_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_15_xor_69_nl = R_7_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_15_xor_70_nl = R_6_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_15_xor_71_nl = R_5_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_15_xor_72_nl = R_4_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_117_rg_addr = {3'b110 , loop_DES_rounds_15_xor_68_nl
      , loop_DES_rounds_15_xor_73_nl , loop_DES_rounds_15_xor_69_nl , loop_DES_rounds_15_xor_70_nl
      , loop_DES_rounds_15_xor_71_nl , loop_DES_rounds_15_xor_72_nl};
  wire[0:0] loop_DES_rounds_15_xor_38_nl;
  wire[0:0] loop_DES_rounds_15_xor_43_nl;
  wire[0:0] loop_DES_rounds_15_xor_39_nl;
  wire[0:0] loop_DES_rounds_15_xor_40_nl;
  wire[0:0] loop_DES_rounds_15_xor_41_nl;
  wire[0:0] loop_DES_rounds_15_xor_42_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_114_rg_addr;
  assign loop_DES_rounds_15_xor_38_nl = R_28_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign loop_DES_rounds_15_xor_43_nl = R_23_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_15_xor_39_nl = R_27_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_15_xor_40_nl = R_26_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_15_xor_41_nl = R_25_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_15_xor_42_nl = R_24_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_114_rg_addr = {3'b001 , loop_DES_rounds_15_xor_38_nl
      , loop_DES_rounds_15_xor_43_nl , loop_DES_rounds_15_xor_39_nl , loop_DES_rounds_15_xor_40_nl
      , loop_DES_rounds_15_xor_41_nl , loop_DES_rounds_15_xor_42_nl};
  wire[0:0] loop_DES_rounds_15_xor_nl;
  wire[0:0] loop_DES_rounds_15_xor_37_nl;
  wire[0:0] loop_DES_rounds_15_xor_33_nl;
  wire[0:0] loop_DES_rounds_15_xor_34_nl;
  wire[0:0] loop_DES_rounds_15_xor_35_nl;
  wire[0:0] loop_DES_rounds_15_xor_36_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_112_rg_addr;
  assign loop_DES_rounds_15_xor_nl = R_0_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign loop_DES_rounds_15_xor_37_nl = R_27_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign loop_DES_rounds_15_xor_33_nl = R_31_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_15_xor_34_nl = R_30_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_15_xor_35_nl = R_29_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_15_xor_36_nl = R_28_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_112_rg_addr = {3'b000 , loop_DES_rounds_15_xor_nl
      , loop_DES_rounds_15_xor_37_nl , loop_DES_rounds_15_xor_33_nl , loop_DES_rounds_15_xor_34_nl
      , loop_DES_rounds_15_xor_35_nl , loop_DES_rounds_15_xor_36_nl};
  wire[0:0] loop_DES_rounds_15_xor_56_nl;
  wire[0:0] loop_DES_rounds_15_xor_61_nl;
  wire[0:0] loop_DES_rounds_15_xor_57_nl;
  wire[0:0] loop_DES_rounds_15_xor_58_nl;
  wire[0:0] loop_DES_rounds_15_xor_59_nl;
  wire[0:0] loop_DES_rounds_15_xor_60_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_113_rg_addr;
  assign loop_DES_rounds_15_xor_56_nl = R_16_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign loop_DES_rounds_15_xor_61_nl = R_11_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_15_xor_57_nl = R_15_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_15_xor_58_nl = R_14_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_15_xor_59_nl = R_13_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign loop_DES_rounds_15_xor_60_nl = R_12_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_113_rg_addr = {3'b100 , loop_DES_rounds_15_xor_56_nl
      , loop_DES_rounds_15_xor_61_nl , loop_DES_rounds_15_xor_57_nl , loop_DES_rounds_15_xor_58_nl
      , loop_DES_rounds_15_xor_59_nl , loop_DES_rounds_15_xor_60_nl};
  wire[0:0] loop_DES_rounds_15_xor_44_nl;
  wire[0:0] loop_DES_rounds_15_xor_49_nl;
  wire[0:0] loop_DES_rounds_15_xor_45_nl;
  wire[0:0] loop_DES_rounds_15_xor_46_nl;
  wire[0:0] loop_DES_rounds_15_xor_47_nl;
  wire[0:0] loop_DES_rounds_15_xor_48_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_116_rg_addr;
  assign loop_DES_rounds_15_xor_44_nl = R_24_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_15_xor_49_nl = R_19_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_15_xor_45_nl = R_23_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_15_xor_46_nl = R_22_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign loop_DES_rounds_15_xor_47_nl = R_21_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_15_xor_48_nl = R_20_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_116_rg_addr = {3'b010 , loop_DES_rounds_15_xor_44_nl
      , loop_DES_rounds_15_xor_49_nl , loop_DES_rounds_15_xor_45_nl , loop_DES_rounds_15_xor_46_nl
      , loop_DES_rounds_15_xor_47_nl , loop_DES_rounds_15_xor_48_nl};
  wire[0:0] loop_DES_rounds_15_xor_62_nl;
  wire[0:0] loop_DES_rounds_15_xor_67_nl;
  wire[0:0] loop_DES_rounds_15_xor_63_nl;
  wire[0:0] loop_DES_rounds_15_xor_64_nl;
  wire[0:0] loop_DES_rounds_15_xor_65_nl;
  wire[0:0] loop_DES_rounds_15_xor_66_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_115_rg_addr;
  assign loop_DES_rounds_15_xor_62_nl = R_12_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_15_xor_67_nl = R_7_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_15_xor_63_nl = R_11_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_15_xor_64_nl = R_10_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_15_xor_65_nl = R_9_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_15_xor_66_nl = R_8_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_115_rg_addr = {3'b101 , loop_DES_rounds_15_xor_62_nl
      , loop_DES_rounds_15_xor_67_nl , loop_DES_rounds_15_xor_63_nl , loop_DES_rounds_15_xor_64_nl
      , loop_DES_rounds_15_xor_65_nl , loop_DES_rounds_15_xor_66_nl};
  wire[0:0] loop_DES_rounds_15_xor_74_nl;
  wire[0:0] loop_DES_rounds_15_xor_79_nl;
  wire[0:0] loop_DES_rounds_15_xor_75_nl;
  wire[0:0] loop_DES_rounds_15_xor_76_nl;
  wire[0:0] loop_DES_rounds_15_xor_77_nl;
  wire[0:0] loop_DES_rounds_15_xor_78_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_119_rg_addr;
  assign loop_DES_rounds_15_xor_74_nl = R_4_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_15_xor_79_nl = R_31_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_15_xor_75_nl = R_3_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_15_xor_76_nl = R_2_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_15_xor_77_nl = R_1_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_15_xor_78_nl = R_0_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_119_rg_addr = {3'b111 , loop_DES_rounds_15_xor_74_nl
      , loop_DES_rounds_15_xor_79_nl , loop_DES_rounds_15_xor_75_nl , loop_DES_rounds_15_xor_76_nl
      , loop_DES_rounds_15_xor_77_nl , loop_DES_rounds_15_xor_78_nl};
  wire[0:0] loop_DES_rounds_16_xor_56_nl;
  wire[0:0] loop_DES_rounds_16_xor_61_nl;
  wire[0:0] loop_DES_rounds_16_xor_57_nl;
  wire[0:0] loop_DES_rounds_16_xor_58_nl;
  wire[0:0] loop_DES_rounds_16_xor_59_nl;
  wire[0:0] loop_DES_rounds_16_xor_60_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_121_rg_addr;
  assign loop_DES_rounds_16_xor_56_nl = R_16_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_16_xor_61_nl = R_11_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_16_xor_57_nl = R_15_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_16_xor_58_nl = R_14_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_16_xor_59_nl = R_13_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_16_xor_60_nl = R_12_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_121_rg_addr = {3'b100 , loop_DES_rounds_16_xor_56_nl
      , loop_DES_rounds_16_xor_61_nl , loop_DES_rounds_16_xor_57_nl , loop_DES_rounds_16_xor_58_nl
      , loop_DES_rounds_16_xor_59_nl , loop_DES_rounds_16_xor_60_nl};
  wire[0:0] loop_DES_rounds_16_xor_nl;
  wire[0:0] loop_DES_rounds_16_xor_37_nl;
  wire[0:0] loop_DES_rounds_16_xor_33_nl;
  wire[0:0] loop_DES_rounds_16_xor_34_nl;
  wire[0:0] loop_DES_rounds_16_xor_35_nl;
  wire[0:0] loop_DES_rounds_16_xor_36_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_120_rg_addr;
  assign loop_DES_rounds_16_xor_nl = R_0_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_16_xor_37_nl = R_27_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_16_xor_33_nl = R_31_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign loop_DES_rounds_16_xor_34_nl = R_30_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign loop_DES_rounds_16_xor_35_nl = R_29_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_16_xor_36_nl = R_28_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_120_rg_addr = {3'b000 , loop_DES_rounds_16_xor_nl
      , loop_DES_rounds_16_xor_37_nl , loop_DES_rounds_16_xor_33_nl , loop_DES_rounds_16_xor_34_nl
      , loop_DES_rounds_16_xor_35_nl , loop_DES_rounds_16_xor_36_nl};
  wire[0:0] loop_DES_rounds_16_xor_44_nl;
  wire[0:0] loop_DES_rounds_16_xor_49_nl;
  wire[0:0] loop_DES_rounds_16_xor_45_nl;
  wire[0:0] loop_DES_rounds_16_xor_46_nl;
  wire[0:0] loop_DES_rounds_16_xor_47_nl;
  wire[0:0] loop_DES_rounds_16_xor_48_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_124_rg_addr;
  assign loop_DES_rounds_16_xor_44_nl = R_24_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_16_xor_49_nl = R_19_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_16_xor_45_nl = R_23_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_16_xor_46_nl = R_22_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_16_xor_47_nl = R_21_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign loop_DES_rounds_16_xor_48_nl = R_20_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_124_rg_addr = {3'b010 , loop_DES_rounds_16_xor_44_nl
      , loop_DES_rounds_16_xor_49_nl , loop_DES_rounds_16_xor_45_nl , loop_DES_rounds_16_xor_46_nl
      , loop_DES_rounds_16_xor_47_nl , loop_DES_rounds_16_xor_48_nl};
  wire[0:0] loop_DES_rounds_16_xor_50_nl;
  wire[0:0] loop_DES_rounds_16_xor_55_nl;
  wire[0:0] loop_DES_rounds_16_xor_51_nl;
  wire[0:0] loop_DES_rounds_16_xor_52_nl;
  wire[0:0] loop_DES_rounds_16_xor_53_nl;
  wire[0:0] loop_DES_rounds_16_xor_54_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_126_rg_addr;
  assign loop_DES_rounds_16_xor_50_nl = R_20_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_16_xor_55_nl = R_15_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign loop_DES_rounds_16_xor_51_nl = R_19_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_16_xor_52_nl = R_18_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_16_xor_53_nl = R_17_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign loop_DES_rounds_16_xor_54_nl = R_16_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_126_rg_addr = {3'b011 , loop_DES_rounds_16_xor_50_nl
      , loop_DES_rounds_16_xor_55_nl , loop_DES_rounds_16_xor_51_nl , loop_DES_rounds_16_xor_52_nl
      , loop_DES_rounds_16_xor_53_nl , loop_DES_rounds_16_xor_54_nl};
  wire[0:0] loop_DES_rounds_16_xor_68_nl;
  wire[0:0] loop_DES_rounds_16_xor_73_nl;
  wire[0:0] loop_DES_rounds_16_xor_69_nl;
  wire[0:0] loop_DES_rounds_16_xor_70_nl;
  wire[0:0] loop_DES_rounds_16_xor_71_nl;
  wire[0:0] loop_DES_rounds_16_xor_72_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_125_rg_addr;
  assign loop_DES_rounds_16_xor_68_nl = R_8_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_16_xor_73_nl = R_3_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_16_xor_69_nl = R_7_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_16_xor_70_nl = R_6_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_16_xor_71_nl = R_5_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_16_xor_72_nl = R_4_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_125_rg_addr = {3'b110 , loop_DES_rounds_16_xor_68_nl
      , loop_DES_rounds_16_xor_73_nl , loop_DES_rounds_16_xor_69_nl , loop_DES_rounds_16_xor_70_nl
      , loop_DES_rounds_16_xor_71_nl , loop_DES_rounds_16_xor_72_nl};
  wire[0:0] loop_DES_rounds_16_xor_38_nl;
  wire[0:0] loop_DES_rounds_16_xor_43_nl;
  wire[0:0] loop_DES_rounds_16_xor_39_nl;
  wire[0:0] loop_DES_rounds_16_xor_40_nl;
  wire[0:0] loop_DES_rounds_16_xor_41_nl;
  wire[0:0] loop_DES_rounds_16_xor_42_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_122_rg_addr;
  assign loop_DES_rounds_16_xor_38_nl = R_28_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_16_xor_43_nl = R_23_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_16_xor_39_nl = R_27_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign loop_DES_rounds_16_xor_40_nl = R_26_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign loop_DES_rounds_16_xor_41_nl = R_25_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_16_xor_42_nl = R_24_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_122_rg_addr = {3'b001 , loop_DES_rounds_16_xor_38_nl
      , loop_DES_rounds_16_xor_43_nl , loop_DES_rounds_16_xor_39_nl , loop_DES_rounds_16_xor_40_nl
      , loop_DES_rounds_16_xor_41_nl , loop_DES_rounds_16_xor_42_nl};
  wire[0:0] loop_DES_rounds_16_xor_74_nl;
  wire[0:0] loop_DES_rounds_16_xor_79_nl;
  wire[0:0] loop_DES_rounds_16_xor_75_nl;
  wire[0:0] loop_DES_rounds_16_xor_76_nl;
  wire[0:0] loop_DES_rounds_16_xor_77_nl;
  wire[0:0] loop_DES_rounds_16_xor_78_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_127_rg_addr;
  assign loop_DES_rounds_16_xor_74_nl = R_4_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_16_xor_79_nl = R_31_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_16_xor_75_nl = R_3_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_16_xor_76_nl = R_2_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_16_xor_77_nl = R_1_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign loop_DES_rounds_16_xor_78_nl = R_0_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_127_rg_addr = {3'b111 , loop_DES_rounds_16_xor_74_nl
      , loop_DES_rounds_16_xor_79_nl , loop_DES_rounds_16_xor_75_nl , loop_DES_rounds_16_xor_76_nl
      , loop_DES_rounds_16_xor_77_nl , loop_DES_rounds_16_xor_78_nl};
  wire[0:0] loop_DES_rounds_16_xor_62_nl;
  wire[0:0] loop_DES_rounds_16_xor_67_nl;
  wire[0:0] loop_DES_rounds_16_xor_63_nl;
  wire[0:0] loop_DES_rounds_16_xor_64_nl;
  wire[0:0] loop_DES_rounds_16_xor_65_nl;
  wire[0:0] loop_DES_rounds_16_xor_66_nl;
  wire [8:0] nl_operator_8_false_1_read_rom_S_rom_map_1_123_rg_addr;
  assign loop_DES_rounds_16_xor_62_nl = R_12_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_16_xor_67_nl = R_7_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_16_xor_63_nl = R_11_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign loop_DES_rounds_16_xor_64_nl = R_10_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_16_xor_65_nl = R_9_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_16_xor_66_nl = R_8_15_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign nl_operator_8_false_1_read_rom_S_rom_map_1_123_rg_addr = {3'b101 , loop_DES_rounds_16_xor_62_nl
      , loop_DES_rounds_16_xor_67_nl , loop_DES_rounds_16_xor_63_nl , loop_DES_rounds_16_xor_64_nl
      , loop_DES_rounds_16_xor_65_nl , loop_DES_rounds_16_xor_66_nl};
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd64)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd64)) key_rsci (
      .dat(key_rsc_dat),
      .idat(key_rsci_idat)
    );
  ccs_out_v1 #(.rscid(32'sd3),
  .width(32'sd64)) return_rsci (
      .idat(nl_return_rsci_idat[63:0]),
      .dat(return_rsc_dat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) input_rsc_triosy_obj (
      .ld(reg_input_rsc_triosy_obj_ld_cse),
      .lz(input_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) key_rsc_triosy_obj (
      .ld(reg_input_rsc_triosy_obj_ld_cse),
      .lz(key_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) return_rsc_triosy_obj (
      .ld(return_rsc_triosy_obj_ld),
      .lz(return_rsc_triosy_lz)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_6_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_6_rg_addr[8:0]),
      .data_out(operator_8_false_1_read_rom_S_rom_map_1_6_itm)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_5_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_5_rg_addr[8:0]),
      .data_out(operator_8_false_1_read_rom_S_rom_map_1_5_itm)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_2_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_2_rg_addr[8:0]),
      .data_out(operator_8_false_1_read_rom_S_rom_map_1_2_itm)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_rg_addr[8:0]),
      .data_out(operator_8_false_1_read_rom_S_rom_map_1_itm)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_1_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_1_rg_addr[8:0]),
      .data_out(operator_8_false_1_read_rom_S_rom_map_1_1_itm)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_4_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_4_rg_addr[8:0]),
      .data_out(operator_8_false_1_read_rom_S_rom_map_1_4_itm)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_3_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_3_rg_addr[8:0]),
      .data_out(operator_8_false_1_read_rom_S_rom_map_1_3_itm)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_7_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_7_rg_addr[8:0]),
      .data_out(operator_8_false_1_read_rom_S_rom_map_1_7_itm)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_14_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_14_rg_addr[8:0]),
      .data_out(operator_8_false_1_read_rom_S_rom_map_1_14_itm)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_13_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_13_rg_addr[8:0]),
      .data_out(operator_8_false_1_read_rom_S_rom_map_1_13_itm)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_10_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_10_rg_addr[8:0]),
      .data_out(operator_8_false_1_read_rom_S_rom_map_1_10_itm)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_8_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_8_rg_addr[8:0]),
      .data_out(operator_8_false_1_read_rom_S_rom_map_1_8_itm)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_9_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_9_rg_addr[8:0]),
      .data_out(operator_8_false_1_read_rom_S_rom_map_1_9_itm)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_12_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_12_rg_addr[8:0]),
      .data_out(operator_8_false_1_read_rom_S_rom_map_1_12_itm)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_11_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_11_rg_addr[8:0]),
      .data_out(operator_8_false_1_read_rom_S_rom_map_1_11_itm)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_15_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_15_rg_addr[8:0]),
      .data_out(operator_8_false_1_read_rom_S_rom_map_1_15_itm)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_22_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_22_rg_addr[8:0]),
      .data_out(s_output_1_19_16_6_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_21_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_21_rg_addr[8:0]),
      .data_out(s_output_1_3_0_55_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_18_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_18_rg_addr[8:0]),
      .data_out(s_output_1_19_16_36_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_16_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_16_rg_addr[8:0]),
      .data_out(s_output_1_19_16_21_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_17_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_17_rg_addr[8:0]),
      .data_out(s_output_1_3_0_25_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_20_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_20_rg_addr[8:0]),
      .data_out(s_output_1_19_16_51_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_19_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_19_rg_addr[8:0]),
      .data_out(s_output_1_3_0_40_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_23_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_23_rg_addr[8:0]),
      .data_out(s_output_1_3_0_10_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_30_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_30_rg_addr[8:0]),
      .data_out(s_output_1_19_16_7_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_29_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_29_rg_addr[8:0]),
      .data_out(s_output_1_3_0_56_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_26_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_26_rg_addr[8:0]),
      .data_out(s_output_1_19_16_37_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_24_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_24_rg_addr[8:0]),
      .data_out(s_output_1_19_16_22_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_25_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_25_rg_addr[8:0]),
      .data_out(s_output_1_3_0_26_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_28_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_28_rg_addr[8:0]),
      .data_out(s_output_1_19_16_52_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_27_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_27_rg_addr[8:0]),
      .data_out(s_output_1_3_0_41_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_31_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_31_rg_addr[8:0]),
      .data_out(s_output_1_3_0_11_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_38_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_38_rg_addr[8:0]),
      .data_out(s_output_1_19_16_8_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_37_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_37_rg_addr[8:0]),
      .data_out(s_output_1_3_0_57_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_34_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_34_rg_addr[8:0]),
      .data_out(s_output_1_19_16_38_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_32_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_32_rg_addr[8:0]),
      .data_out(s_output_1_19_16_23_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_33_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_33_rg_addr[8:0]),
      .data_out(s_output_1_3_0_27_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_36_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_36_rg_addr[8:0]),
      .data_out(s_output_1_19_16_53_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_35_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_35_rg_addr[8:0]),
      .data_out(s_output_1_3_0_42_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_39_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_39_rg_addr[8:0]),
      .data_out(s_output_1_3_0_12_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_46_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_46_rg_addr[8:0]),
      .data_out(s_output_1_19_16_9_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_45_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_45_rg_addr[8:0]),
      .data_out(s_output_1_3_0_58_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_42_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_42_rg_addr[8:0]),
      .data_out(s_output_1_19_16_39_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_40_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_40_rg_addr[8:0]),
      .data_out(s_output_1_19_16_24_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_41_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_41_rg_addr[8:0]),
      .data_out(s_output_1_3_0_28_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_44_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_44_rg_addr[8:0]),
      .data_out(s_output_1_19_16_54_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_43_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_43_rg_addr[8:0]),
      .data_out(s_output_1_3_0_43_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_47_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_47_rg_addr[8:0]),
      .data_out(s_output_1_3_0_13_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_54_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_54_rg_addr[8:0]),
      .data_out(s_output_1_19_16_10_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_53_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_53_rg_addr[8:0]),
      .data_out(s_output_1_3_0_59_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_50_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_50_rg_addr[8:0]),
      .data_out(s_output_1_19_16_40_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_48_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_48_rg_addr[8:0]),
      .data_out(s_output_1_19_16_25_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_49_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_49_rg_addr[8:0]),
      .data_out(s_output_1_3_0_29_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_52_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_52_rg_addr[8:0]),
      .data_out(s_output_1_19_16_55_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_51_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_51_rg_addr[8:0]),
      .data_out(s_output_1_3_0_44_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_55_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_55_rg_addr[8:0]),
      .data_out(s_output_1_3_0_14_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_62_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_62_rg_addr[8:0]),
      .data_out(s_output_1_19_16_11_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_61_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_61_rg_addr[8:0]),
      .data_out(s_output_1_3_0_60_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_58_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_58_rg_addr[8:0]),
      .data_out(s_output_1_19_16_41_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_56_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_56_rg_addr[8:0]),
      .data_out(s_output_1_19_16_26_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_57_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_57_rg_addr[8:0]),
      .data_out(s_output_1_3_0_30_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_60_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_60_rg_addr[8:0]),
      .data_out(s_output_1_19_16_56_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_59_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_59_rg_addr[8:0]),
      .data_out(s_output_1_3_0_45_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_63_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_63_rg_addr[8:0]),
      .data_out(s_output_1_3_0_15_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_70_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_70_rg_addr[8:0]),
      .data_out(s_output_1_19_16_12_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_69_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_69_rg_addr[8:0]),
      .data_out(s_output_1_3_0_61_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_66_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_66_rg_addr[8:0]),
      .data_out(s_output_1_19_16_42_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_64_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_64_rg_addr[8:0]),
      .data_out(s_output_1_19_16_27_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_65_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_65_rg_addr[8:0]),
      .data_out(s_output_1_3_0_31_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_68_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_68_rg_addr[8:0]),
      .data_out(s_output_1_19_16_57_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_67_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_67_rg_addr[8:0]),
      .data_out(s_output_1_3_0_46_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_71_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_71_rg_addr[8:0]),
      .data_out(s_output_1_3_0_16_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_78_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_78_rg_addr[8:0]),
      .data_out(s_output_1_19_16_13_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_77_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_77_rg_addr[8:0]),
      .data_out(s_output_1_3_0_62_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_74_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_74_rg_addr[8:0]),
      .data_out(s_output_1_19_16_43_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_72_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_72_rg_addr[8:0]),
      .data_out(s_output_1_19_16_28_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_73_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_73_rg_addr[8:0]),
      .data_out(s_output_1_3_0_32_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_76_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_76_rg_addr[8:0]),
      .data_out(s_output_1_19_16_58_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_75_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_75_rg_addr[8:0]),
      .data_out(s_output_1_3_0_47_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_79_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_79_rg_addr[8:0]),
      .data_out(s_output_1_3_0_17_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_86_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_86_rg_addr[8:0]),
      .data_out(s_output_1_19_16_14_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_85_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_85_rg_addr[8:0]),
      .data_out(s_output_1_3_0_63_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_82_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_82_rg_addr[8:0]),
      .data_out(s_output_1_19_16_44_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_80_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_80_rg_addr[8:0]),
      .data_out(s_output_1_19_16_29_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_81_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_81_rg_addr[8:0]),
      .data_out(s_output_1_3_0_33_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_84_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_84_rg_addr[8:0]),
      .data_out(s_output_1_19_16_59_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_83_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_83_rg_addr[8:0]),
      .data_out(s_output_1_3_0_48_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_87_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_87_rg_addr[8:0]),
      .data_out(s_output_1_3_0_18_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_94_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_94_rg_addr[8:0]),
      .data_out(s_output_1_19_16_15_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_93_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_93_rg_addr[8:0]),
      .data_out(s_output_1_3_0_64_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_90_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_90_rg_addr[8:0]),
      .data_out(s_output_1_19_16_45_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_88_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_88_rg_addr[8:0]),
      .data_out(s_output_1_19_16_30_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_89_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_89_rg_addr[8:0]),
      .data_out(s_output_1_3_0_34_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_92_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_92_rg_addr[8:0]),
      .data_out(s_output_1_19_16_60_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_91_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_91_rg_addr[8:0]),
      .data_out(s_output_1_3_0_49_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_95_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_95_rg_addr[8:0]),
      .data_out(s_output_1_3_0_19_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_102_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_102_rg_addr[8:0]),
      .data_out(s_output_1_19_16_16_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_101_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_101_rg_addr[8:0]),
      .data_out(s_output_1_3_0_65_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_98_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_98_rg_addr[8:0]),
      .data_out(s_output_1_19_16_46_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_96_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_96_rg_addr[8:0]),
      .data_out(s_output_1_19_16_31_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_97_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_97_rg_addr[8:0]),
      .data_out(s_output_1_3_0_35_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_100_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_100_rg_addr[8:0]),
      .data_out(s_output_1_19_16_61_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_99_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_99_rg_addr[8:0]),
      .data_out(s_output_1_3_0_50_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_103_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_103_rg_addr[8:0]),
      .data_out(s_output_1_3_0_20_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_110_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_110_rg_addr[8:0]),
      .data_out(s_output_1_19_16_17_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_109_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_109_rg_addr[8:0]),
      .data_out(s_output_1_3_0_66_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_106_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_106_rg_addr[8:0]),
      .data_out(s_output_1_19_16_47_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_104_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_104_rg_addr[8:0]),
      .data_out(s_output_1_19_16_32_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_105_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_105_rg_addr[8:0]),
      .data_out(s_output_1_3_0_36_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_108_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_108_rg_addr[8:0]),
      .data_out(s_output_1_19_16_62_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_107_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_107_rg_addr[8:0]),
      .data_out(s_output_1_3_0_51_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_111_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_111_rg_addr[8:0]),
      .data_out(s_output_1_3_0_21_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_118_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_118_rg_addr[8:0]),
      .data_out(s_output_1_19_16_18_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_117_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_117_rg_addr[8:0]),
      .data_out(s_output_1_3_0_67_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_114_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_114_rg_addr[8:0]),
      .data_out(s_output_1_19_16_48_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_112_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_112_rg_addr[8:0]),
      .data_out(s_output_1_19_16_33_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_113_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_113_rg_addr[8:0]),
      .data_out(s_output_1_3_0_37_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_116_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_116_rg_addr[8:0]),
      .data_out(s_output_1_19_16_63_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_115_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_115_rg_addr[8:0]),
      .data_out(s_output_1_3_0_52_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_119_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_119_rg_addr[8:0]),
      .data_out(s_output_1_3_0_22_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_121_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_121_rg_addr[8:0]),
      .data_out(s_output_1_3_0_5_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_120_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_120_rg_addr[8:0]),
      .data_out(s_output_1_19_16_1_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_124_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_124_rg_addr[8:0]),
      .data_out(s_output_1_19_16_3_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_126_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_126_rg_addr[8:0]),
      .data_out(s_output_1_19_16_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_125_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_125_rg_addr[8:0]),
      .data_out(s_output_1_3_0_7_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_122_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_122_rg_addr[8:0]),
      .data_out(s_output_1_19_16_2_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_127_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_127_rg_addr[8:0]),
      .data_out(s_output_1_3_0_sva_1)
    );
  des_checkmgc_rom_12_512_4_1  operator_8_false_1_read_rom_S_rom_map_1_123_rg (
      .addr(nl_operator_8_false_1_read_rom_S_rom_map_1_123_rg_addr[8:0]),
      .data_out(s_output_1_3_0_6_sva_1)
    );
  des_check_core_core_fsm des_check_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output)
    );
  always @(posedge clk) begin
    if ( fsm_output[0] ) begin
      key_io_read_key_rsc_cse_63_1_sva <= key_rsci_idat[63:1];
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_31 <= R_28_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_32 <= R_3_14_sva ^ (s_output_1_3_0_6_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_30 <= R_28_14_sva ^ (s_output_1_3_0_6_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_33 <= R_3_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_29 <= R_20_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_34 <= R_11_14_sva ^ (s_output_1_3_0_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_28 <= R_20_14_sva ^ (s_output_1_3_0_7_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_35 <= R_11_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_27 <= R_12_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_36 <= R_19_14_sva ^ (s_output_1_19_16_2_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_26 <= R_12_14_sva ^ (s_output_1_19_16_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_37 <= R_19_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_25 <= R_4_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_38 <= R_27_14_sva ^ (s_output_1_3_0_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_24 <= R_4_14_sva ^ (s_output_1_19_16_2_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_39 <= R_27_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_23 <= R_29_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_40 <= R_2_14_sva ^ (s_output_1_19_16_3_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_22 <= R_29_14_sva ^ (s_output_1_3_0_5_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_41 <= R_2_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_21 <= R_21_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_42 <= R_10_14_sva ^ (s_output_1_3_0_7_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_20 <= R_21_14_sva ^ (s_output_1_3_0_6_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_43 <= R_10_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_19 <= R_13_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_44 <= R_18_14_sva ^ (s_output_1_3_0_5_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_18 <= R_13_14_sva ^ (s_output_1_3_0_6_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_45 <= R_18_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_17 <= R_5_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_46 <= R_26_14_sva ^ (s_output_1_19_16_3_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_16 <= R_5_14_sva ^ (s_output_1_3_0_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_47 <= R_26_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_15 <= R_30_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_48 <= R_1_14_sva ^ (s_output_1_19_16_1_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_14 <= R_30_14_sva ^ (s_output_1_19_16_2_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_49 <= R_1_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_13 <= R_22_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_50 <= R_9_14_sva ^ (s_output_1_19_16_1_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_12 <= R_22_14_sva ^ (s_output_1_19_16_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_51 <= R_9_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_11 <= R_14_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_52 <= R_17_14_sva ^ (s_output_1_3_0_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_10 <= R_14_14_sva ^ (s_output_1_19_16_2_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_53 <= R_17_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_9 <= R_6_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_54 <= R_25_14_sva ^ (s_output_1_3_0_7_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_8 <= R_6_14_sva ^ (s_output_1_19_16_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_55 <= R_25_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_7 <= R_31_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_56 <= R_0_14_sva ^ (s_output_1_3_0_7_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_6 <= R_31_14_sva ^ (s_output_1_19_16_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_57 <= R_0_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_5 <= R_23_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_58 <= R_8_14_sva ^ (s_output_1_19_16_3_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_4 <= R_23_14_sva ^ (s_output_1_19_16_1_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_59 <= R_8_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_3 <= R_15_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_60 <= R_16_14_sva ^ (s_output_1_19_16_3_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_2 <= R_15_14_sva ^ (s_output_1_19_16_1_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_61 <= R_16_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_1 <= R_7_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_62 <= R_24_14_sva ^ (s_output_1_3_0_5_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_0 <= R_7_14_sva ^ (s_output_1_3_0_5_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[15] ) begin
      return_rsci_idat_63 <= R_24_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[0] ) begin
      input_sva <= input_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_input_rsc_triosy_obj_ld_cse <= 1'b0;
      return_rsc_triosy_obj_ld <= 1'b0;
    end
    else begin
      reg_input_rsc_triosy_obj_ld_cse <= fsm_output[0];
      return_rsc_triosy_obj_ld <= fsm_output[15];
    end
  end
  always @(posedge clk) begin
    s_output_1_19_16_4_sva <= operator_8_false_1_read_rom_S_rom_map_1_6_itm;
    s_output_1_3_0_53_sva <= operator_8_false_1_read_rom_S_rom_map_1_5_itm;
    s_output_1_19_16_34_sva <= operator_8_false_1_read_rom_S_rom_map_1_2_itm;
    s_output_1_19_16_19_sva <= operator_8_false_1_read_rom_S_rom_map_1_itm;
    s_output_1_3_0_23_sva <= operator_8_false_1_read_rom_S_rom_map_1_1_itm;
    s_output_1_19_16_49_sva <= operator_8_false_1_read_rom_S_rom_map_1_4_itm;
    s_output_1_3_0_38_sva <= operator_8_false_1_read_rom_S_rom_map_1_3_itm;
    s_output_1_3_0_8_sva <= operator_8_false_1_read_rom_S_rom_map_1_7_itm;
    R_31_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_32_nl, loop_DES_rounds_2_xor_32_nl,
        fsm_output[2]);
    R_0_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_31_nl, loop_DES_rounds_2_xor_31_nl,
        fsm_output[2]);
    R_30_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_30_nl, loop_DES_rounds_2_xor_30_nl,
        fsm_output[2]);
    R_1_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_29_nl, loop_DES_rounds_2_xor_29_nl,
        fsm_output[2]);
    R_29_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_28_nl, loop_DES_rounds_2_xor_28_nl,
        fsm_output[2]);
    R_2_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_27_nl, loop_DES_rounds_2_xor_27_nl,
        fsm_output[2]);
    R_28_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_26_nl, loop_DES_rounds_2_xor_26_nl,
        fsm_output[2]);
    R_3_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_25_nl, loop_DES_rounds_2_xor_25_nl,
        fsm_output[2]);
    R_27_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_24_nl, loop_DES_rounds_2_xor_24_nl,
        fsm_output[2]);
    R_4_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_23_nl, loop_DES_rounds_2_xor_23_nl,
        fsm_output[2]);
    R_26_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_22_nl, loop_DES_rounds_2_xor_22_nl,
        fsm_output[2]);
    R_5_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_21_nl, loop_DES_rounds_2_xor_21_nl,
        fsm_output[2]);
    R_25_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_20_nl, loop_DES_rounds_2_xor_20_nl,
        fsm_output[2]);
    R_6_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_19_nl, loop_DES_rounds_2_xor_19_nl,
        fsm_output[2]);
    R_24_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_18_nl, loop_DES_rounds_2_xor_18_nl,
        fsm_output[2]);
    R_7_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_17_nl, loop_DES_rounds_2_xor_17_nl,
        fsm_output[2]);
    R_23_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_16_nl, loop_DES_rounds_2_xor_16_nl,
        fsm_output[2]);
    R_8_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_15_nl, loop_DES_rounds_2_xor_15_nl,
        fsm_output[2]);
    R_22_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_14_nl, loop_DES_rounds_2_xor_14_nl,
        fsm_output[2]);
    R_9_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_13_nl, loop_DES_rounds_2_xor_13_nl,
        fsm_output[2]);
    R_21_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_12_nl, loop_DES_rounds_2_xor_12_nl,
        fsm_output[2]);
    R_10_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_11_nl, loop_DES_rounds_2_xor_11_nl,
        fsm_output[2]);
    R_20_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_10_nl, loop_DES_rounds_2_xor_10_nl,
        fsm_output[2]);
    R_11_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_9_nl, loop_DES_rounds_2_xor_9_nl,
        fsm_output[2]);
    R_19_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_8_nl, loop_DES_rounds_2_xor_8_nl,
        fsm_output[2]);
    R_12_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_7_nl, loop_DES_rounds_2_xor_7_nl,
        fsm_output[2]);
    R_18_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_6_nl, loop_DES_rounds_2_xor_6_nl,
        fsm_output[2]);
    R_13_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_5_nl, loop_DES_rounds_2_xor_5_nl,
        fsm_output[2]);
    R_17_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_4_nl, loop_DES_rounds_2_xor_4_nl,
        fsm_output[2]);
    R_14_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_3_nl, loop_DES_rounds_2_xor_3_nl,
        fsm_output[2]);
    R_16_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_2_nl, loop_DES_rounds_2_xor_2_nl,
        fsm_output[2]);
    R_15_1_sva <= MUX_s_1_2_2(loop_DES_rounds_1_xor_1_nl, loop_DES_rounds_2_xor_1_nl,
        fsm_output[2]);
    s_output_1_19_16_5_sva <= operator_8_false_1_read_rom_S_rom_map_1_14_itm;
    s_output_1_3_0_54_sva <= operator_8_false_1_read_rom_S_rom_map_1_13_itm;
    s_output_1_19_16_35_sva <= operator_8_false_1_read_rom_S_rom_map_1_10_itm;
    s_output_1_19_16_20_sva <= operator_8_false_1_read_rom_S_rom_map_1_8_itm;
    s_output_1_3_0_24_sva <= operator_8_false_1_read_rom_S_rom_map_1_9_itm;
    s_output_1_19_16_50_sva <= operator_8_false_1_read_rom_S_rom_map_1_12_itm;
    s_output_1_3_0_39_sva <= operator_8_false_1_read_rom_S_rom_map_1_11_itm;
    s_output_1_3_0_9_sva <= operator_8_false_1_read_rom_S_rom_map_1_15_itm;
    R_24_15_sva <= R_24_13_sva ^ (s_output_1_3_0_37_sva_1[3]);
    R_7_15_sva <= R_7_13_sva ^ (s_output_1_3_0_37_sva_1[1]);
    R_16_15_sva <= R_16_13_sva ^ (s_output_1_19_16_63_sva_1[2]);
    R_15_15_sva <= R_15_13_sva ^ (s_output_1_19_16_33_sva_1[2]);
    R_8_15_sva <= R_8_13_sva ^ (s_output_1_19_16_63_sva_1[3]);
    R_23_15_sva <= R_23_13_sva ^ (s_output_1_19_16_33_sva_1[3]);
    R_0_15_sva <= R_0_13_sva ^ (s_output_1_3_0_67_sva_1[3]);
    R_31_15_sva <= R_31_13_sva ^ (s_output_1_19_16_18_sva_1[0]);
    R_25_15_sva <= R_25_13_sva ^ (s_output_1_3_0_67_sva_1[0]);
    R_6_15_sva <= R_6_13_sva ^ (s_output_1_19_16_18_sva_1[3]);
    R_17_15_sva <= R_17_13_sva ^ (s_output_1_3_0_22_sva_1[1]);
    R_14_15_sva <= R_14_13_sva ^ (s_output_1_19_16_48_sva_1[0]);
    R_9_15_sva <= R_9_13_sva ^ (s_output_1_19_16_33_sva_1[1]);
    R_22_15_sva <= R_22_13_sva ^ (s_output_1_19_16_18_sva_1[1]);
    R_1_15_sva <= R_1_13_sva ^ (s_output_1_19_16_33_sva_1[0]);
    R_30_15_sva <= R_30_13_sva ^ (s_output_1_19_16_48_sva_1[1]);
    R_26_15_sva <= R_26_13_sva ^ (s_output_1_19_16_63_sva_1[0]);
    R_5_15_sva <= R_5_13_sva ^ (s_output_1_3_0_22_sva_1[2]);
    R_18_15_sva <= R_18_13_sva ^ (s_output_1_3_0_37_sva_1[2]);
    R_13_15_sva <= R_13_13_sva ^ (s_output_1_3_0_52_sva_1[0]);
    R_10_15_sva <= R_10_13_sva ^ (s_output_1_3_0_67_sva_1[1]);
    R_21_15_sva <= R_21_13_sva ^ (s_output_1_3_0_52_sva_1[1]);
    R_2_15_sva <= R_2_13_sva ^ (s_output_1_19_16_63_sva_1[1]);
    R_29_15_sva <= R_29_13_sva ^ (s_output_1_3_0_37_sva_1[0]);
    R_27_15_sva <= R_27_13_sva ^ (s_output_1_3_0_22_sva_1[3]);
    R_4_15_sva <= R_4_13_sva ^ (s_output_1_19_16_48_sva_1[2]);
    R_19_15_sva <= R_19_13_sva ^ (s_output_1_19_16_48_sva_1[3]);
    R_12_15_sva <= R_12_13_sva ^ (s_output_1_19_16_18_sva_1[2]);
    R_11_15_sva <= R_11_13_sva ^ (s_output_1_3_0_22_sva_1[0]);
    R_20_15_sva <= R_20_13_sva ^ (s_output_1_3_0_67_sva_1[2]);
    R_3_15_sva <= R_3_13_sva ^ (s_output_1_3_0_52_sva_1[2]);
    R_28_15_sva <= R_28_13_sva ^ (s_output_1_3_0_52_sva_1[3]);
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_31_3_sva <= R_31_1_sva ^ (s_output_1_19_16_6_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_0_3_sva <= R_0_1_sva ^ (s_output_1_3_0_55_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_30_3_sva <= R_30_1_sva ^ (s_output_1_19_16_36_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_1_3_sva <= R_1_1_sva ^ (s_output_1_19_16_21_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_29_3_sva <= R_29_1_sva ^ (s_output_1_3_0_25_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_2_3_sva <= R_2_1_sva ^ (s_output_1_19_16_51_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_28_3_sva <= R_28_1_sva ^ (s_output_1_3_0_40_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_3_3_sva <= R_3_1_sva ^ (s_output_1_3_0_40_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_27_3_sva <= R_27_1_sva ^ (s_output_1_3_0_10_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_4_3_sva <= R_4_1_sva ^ (s_output_1_19_16_36_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_26_3_sva <= R_26_1_sva ^ (s_output_1_19_16_51_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_5_3_sva <= R_5_1_sva ^ (s_output_1_3_0_10_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_25_3_sva <= R_25_1_sva ^ (s_output_1_3_0_55_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_6_3_sva <= R_6_1_sva ^ (s_output_1_19_16_6_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_24_3_sva <= R_24_1_sva ^ (s_output_1_3_0_25_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_7_3_sva <= R_7_1_sva ^ (s_output_1_3_0_25_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_23_3_sva <= R_23_1_sva ^ (s_output_1_19_16_21_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_8_3_sva <= R_8_1_sva ^ (s_output_1_19_16_51_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_22_3_sva <= R_22_1_sva ^ (s_output_1_19_16_6_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_9_3_sva <= R_9_1_sva ^ (s_output_1_19_16_21_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_21_3_sva <= R_21_1_sva ^ (s_output_1_3_0_40_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_10_3_sva <= R_10_1_sva ^ (s_output_1_3_0_55_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_20_3_sva <= R_20_1_sva ^ (s_output_1_3_0_55_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_11_3_sva <= R_11_1_sva ^ (s_output_1_3_0_10_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_19_3_sva <= R_19_1_sva ^ (s_output_1_19_16_36_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_12_3_sva <= R_12_1_sva ^ (s_output_1_19_16_6_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_18_3_sva <= R_18_1_sva ^ (s_output_1_3_0_25_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_13_3_sva <= R_13_1_sva ^ (s_output_1_3_0_40_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_17_3_sva <= R_17_1_sva ^ (s_output_1_3_0_10_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_14_3_sva <= R_14_1_sva ^ (s_output_1_19_16_36_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_16_3_sva <= R_16_1_sva ^ (s_output_1_19_16_51_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[2] ) begin
      R_15_3_sva <= R_15_1_sva ^ (s_output_1_19_16_21_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_31_4_sva <= R_31_1_sva ^ (s_output_1_19_16_7_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_0_4_sva <= R_0_1_sva ^ (s_output_1_3_0_56_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_30_4_sva <= R_30_1_sva ^ (s_output_1_19_16_37_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_1_4_sva <= R_1_1_sva ^ (s_output_1_19_16_22_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_29_4_sva <= R_29_1_sva ^ (s_output_1_3_0_26_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_2_4_sva <= R_2_1_sva ^ (s_output_1_19_16_52_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_28_4_sva <= R_28_1_sva ^ (s_output_1_3_0_41_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_3_4_sva <= R_3_1_sva ^ (s_output_1_3_0_41_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_27_4_sva <= R_27_1_sva ^ (s_output_1_3_0_11_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_4_4_sva <= R_4_1_sva ^ (s_output_1_19_16_37_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_26_4_sva <= R_26_1_sva ^ (s_output_1_19_16_52_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_5_4_sva <= R_5_1_sva ^ (s_output_1_3_0_11_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_25_4_sva <= R_25_1_sva ^ (s_output_1_3_0_56_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_6_4_sva <= R_6_1_sva ^ (s_output_1_19_16_7_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_24_4_sva <= R_24_1_sva ^ (s_output_1_3_0_26_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_7_4_sva <= R_7_1_sva ^ (s_output_1_3_0_26_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_23_4_sva <= R_23_1_sva ^ (s_output_1_19_16_22_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_8_4_sva <= R_8_1_sva ^ (s_output_1_19_16_52_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_22_4_sva <= R_22_1_sva ^ (s_output_1_19_16_7_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_9_4_sva <= R_9_1_sva ^ (s_output_1_19_16_22_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_21_4_sva <= R_21_1_sva ^ (s_output_1_3_0_41_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_10_4_sva <= R_10_1_sva ^ (s_output_1_3_0_56_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_20_4_sva <= R_20_1_sva ^ (s_output_1_3_0_56_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_11_4_sva <= R_11_1_sva ^ (s_output_1_3_0_11_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_19_4_sva <= R_19_1_sva ^ (s_output_1_19_16_37_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_12_4_sva <= R_12_1_sva ^ (s_output_1_19_16_7_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_18_4_sva <= R_18_1_sva ^ (s_output_1_3_0_26_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_13_4_sva <= R_13_1_sva ^ (s_output_1_3_0_41_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_17_4_sva <= R_17_1_sva ^ (s_output_1_3_0_11_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_14_4_sva <= R_14_1_sva ^ (s_output_1_19_16_37_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_16_4_sva <= R_16_1_sva ^ (s_output_1_19_16_52_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[3] ) begin
      R_15_4_sva <= R_15_1_sva ^ (s_output_1_19_16_22_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_31_5_sva <= R_31_3_sva ^ (s_output_1_19_16_8_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_0_5_sva <= R_0_3_sva ^ (s_output_1_3_0_57_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_30_5_sva <= R_30_3_sva ^ (s_output_1_19_16_38_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_1_5_sva <= R_1_3_sva ^ (s_output_1_19_16_23_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_29_5_sva <= R_29_3_sva ^ (s_output_1_3_0_27_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_2_5_sva <= R_2_3_sva ^ (s_output_1_19_16_53_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_28_5_sva <= R_28_3_sva ^ (s_output_1_3_0_42_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_3_5_sva <= R_3_3_sva ^ (s_output_1_3_0_42_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_27_5_sva <= R_27_3_sva ^ (s_output_1_3_0_12_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_4_5_sva <= R_4_3_sva ^ (s_output_1_19_16_38_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_26_5_sva <= R_26_3_sva ^ (s_output_1_19_16_53_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_5_5_sva <= R_5_3_sva ^ (s_output_1_3_0_12_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_25_5_sva <= R_25_3_sva ^ (s_output_1_3_0_57_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_6_5_sva <= R_6_3_sva ^ (s_output_1_19_16_8_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_24_5_sva <= R_24_3_sva ^ (s_output_1_3_0_27_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_7_5_sva <= R_7_3_sva ^ (s_output_1_3_0_27_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_23_5_sva <= R_23_3_sva ^ (s_output_1_19_16_23_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_8_5_sva <= R_8_3_sva ^ (s_output_1_19_16_53_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_22_5_sva <= R_22_3_sva ^ (s_output_1_19_16_8_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_9_5_sva <= R_9_3_sva ^ (s_output_1_19_16_23_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_21_5_sva <= R_21_3_sva ^ (s_output_1_3_0_42_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_10_5_sva <= R_10_3_sva ^ (s_output_1_3_0_57_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_20_5_sva <= R_20_3_sva ^ (s_output_1_3_0_57_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_11_5_sva <= R_11_3_sva ^ (s_output_1_3_0_12_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_19_5_sva <= R_19_3_sva ^ (s_output_1_19_16_38_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_12_5_sva <= R_12_3_sva ^ (s_output_1_19_16_8_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_18_5_sva <= R_18_3_sva ^ (s_output_1_3_0_27_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_13_5_sva <= R_13_3_sva ^ (s_output_1_3_0_42_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_17_5_sva <= R_17_3_sva ^ (s_output_1_3_0_12_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_14_5_sva <= R_14_3_sva ^ (s_output_1_19_16_38_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_16_5_sva <= R_16_3_sva ^ (s_output_1_19_16_53_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[4] ) begin
      R_15_5_sva <= R_15_3_sva ^ (s_output_1_19_16_23_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_31_6_sva <= R_31_4_sva ^ (s_output_1_19_16_9_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_0_6_sva <= R_0_4_sva ^ (s_output_1_3_0_58_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_30_6_sva <= R_30_4_sva ^ (s_output_1_19_16_39_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_1_6_sva <= R_1_4_sva ^ (s_output_1_19_16_24_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_29_6_sva <= R_29_4_sva ^ (s_output_1_3_0_28_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_2_6_sva <= R_2_4_sva ^ (s_output_1_19_16_54_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_28_6_sva <= R_28_4_sva ^ (s_output_1_3_0_43_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_3_6_sva <= R_3_4_sva ^ (s_output_1_3_0_43_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_27_6_sva <= R_27_4_sva ^ (s_output_1_3_0_13_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_4_6_sva <= R_4_4_sva ^ (s_output_1_19_16_39_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_26_6_sva <= R_26_4_sva ^ (s_output_1_19_16_54_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_5_6_sva <= R_5_4_sva ^ (s_output_1_3_0_13_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_25_6_sva <= R_25_4_sva ^ (s_output_1_3_0_58_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_6_6_sva <= R_6_4_sva ^ (s_output_1_19_16_9_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_24_6_sva <= R_24_4_sva ^ (s_output_1_3_0_28_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_7_6_sva <= R_7_4_sva ^ (s_output_1_3_0_28_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_23_6_sva <= R_23_4_sva ^ (s_output_1_19_16_24_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_8_6_sva <= R_8_4_sva ^ (s_output_1_19_16_54_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_22_6_sva <= R_22_4_sva ^ (s_output_1_19_16_9_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_9_6_sva <= R_9_4_sva ^ (s_output_1_19_16_24_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_21_6_sva <= R_21_4_sva ^ (s_output_1_3_0_43_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_10_6_sva <= R_10_4_sva ^ (s_output_1_3_0_58_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_20_6_sva <= R_20_4_sva ^ (s_output_1_3_0_58_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_11_6_sva <= R_11_4_sva ^ (s_output_1_3_0_13_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_19_6_sva <= R_19_4_sva ^ (s_output_1_19_16_39_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_12_6_sva <= R_12_4_sva ^ (s_output_1_19_16_9_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_18_6_sva <= R_18_4_sva ^ (s_output_1_3_0_28_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_13_6_sva <= R_13_4_sva ^ (s_output_1_3_0_43_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_17_6_sva <= R_17_4_sva ^ (s_output_1_3_0_13_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_14_6_sva <= R_14_4_sva ^ (s_output_1_19_16_39_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_16_6_sva <= R_16_4_sva ^ (s_output_1_19_16_54_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      R_15_6_sva <= R_15_4_sva ^ (s_output_1_19_16_24_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_31_7_sva <= R_31_5_sva ^ (s_output_1_19_16_10_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_0_7_sva <= R_0_5_sva ^ (s_output_1_3_0_59_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_30_7_sva <= R_30_5_sva ^ (s_output_1_19_16_40_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_1_7_sva <= R_1_5_sva ^ (s_output_1_19_16_25_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_29_7_sva <= R_29_5_sva ^ (s_output_1_3_0_29_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_2_7_sva <= R_2_5_sva ^ (s_output_1_19_16_55_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_28_7_sva <= R_28_5_sva ^ (s_output_1_3_0_44_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_3_7_sva <= R_3_5_sva ^ (s_output_1_3_0_44_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_27_7_sva <= R_27_5_sva ^ (s_output_1_3_0_14_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_4_7_sva <= R_4_5_sva ^ (s_output_1_19_16_40_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_26_7_sva <= R_26_5_sva ^ (s_output_1_19_16_55_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_5_7_sva <= R_5_5_sva ^ (s_output_1_3_0_14_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_25_7_sva <= R_25_5_sva ^ (s_output_1_3_0_59_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_6_7_sva <= R_6_5_sva ^ (s_output_1_19_16_10_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_24_7_sva <= R_24_5_sva ^ (s_output_1_3_0_29_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_7_7_sva <= R_7_5_sva ^ (s_output_1_3_0_29_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_23_7_sva <= R_23_5_sva ^ (s_output_1_19_16_25_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_8_7_sva <= R_8_5_sva ^ (s_output_1_19_16_55_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_22_7_sva <= R_22_5_sva ^ (s_output_1_19_16_10_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_9_7_sva <= R_9_5_sva ^ (s_output_1_19_16_25_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_21_7_sva <= R_21_5_sva ^ (s_output_1_3_0_44_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_10_7_sva <= R_10_5_sva ^ (s_output_1_3_0_59_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_20_7_sva <= R_20_5_sva ^ (s_output_1_3_0_59_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_11_7_sva <= R_11_5_sva ^ (s_output_1_3_0_14_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_19_7_sva <= R_19_5_sva ^ (s_output_1_19_16_40_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_12_7_sva <= R_12_5_sva ^ (s_output_1_19_16_10_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_18_7_sva <= R_18_5_sva ^ (s_output_1_3_0_29_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_13_7_sva <= R_13_5_sva ^ (s_output_1_3_0_44_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_17_7_sva <= R_17_5_sva ^ (s_output_1_3_0_14_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_14_7_sva <= R_14_5_sva ^ (s_output_1_19_16_40_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_16_7_sva <= R_16_5_sva ^ (s_output_1_19_16_55_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[6] ) begin
      R_15_7_sva <= R_15_5_sva ^ (s_output_1_19_16_25_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_31_8_sva <= R_31_6_sva ^ (s_output_1_19_16_11_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_0_8_sva <= R_0_6_sva ^ (s_output_1_3_0_60_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_30_8_sva <= R_30_6_sva ^ (s_output_1_19_16_41_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_1_8_sva <= R_1_6_sva ^ (s_output_1_19_16_26_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_29_8_sva <= R_29_6_sva ^ (s_output_1_3_0_30_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_2_8_sva <= R_2_6_sva ^ (s_output_1_19_16_56_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_28_8_sva <= R_28_6_sva ^ (s_output_1_3_0_45_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_3_8_sva <= R_3_6_sva ^ (s_output_1_3_0_45_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_27_8_sva <= R_27_6_sva ^ (s_output_1_3_0_15_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_4_8_sva <= R_4_6_sva ^ (s_output_1_19_16_41_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_26_8_sva <= R_26_6_sva ^ (s_output_1_19_16_56_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_5_8_sva <= R_5_6_sva ^ (s_output_1_3_0_15_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_25_8_sva <= R_25_6_sva ^ (s_output_1_3_0_60_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_6_8_sva <= R_6_6_sva ^ (s_output_1_19_16_11_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_24_8_sva <= R_24_6_sva ^ (s_output_1_3_0_30_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_7_8_sva <= R_7_6_sva ^ (s_output_1_3_0_30_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_23_8_sva <= R_23_6_sva ^ (s_output_1_19_16_26_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_8_8_sva <= R_8_6_sva ^ (s_output_1_19_16_56_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_22_8_sva <= R_22_6_sva ^ (s_output_1_19_16_11_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_9_8_sva <= R_9_6_sva ^ (s_output_1_19_16_26_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_21_8_sva <= R_21_6_sva ^ (s_output_1_3_0_45_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_10_8_sva <= R_10_6_sva ^ (s_output_1_3_0_60_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_20_8_sva <= R_20_6_sva ^ (s_output_1_3_0_60_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_11_8_sva <= R_11_6_sva ^ (s_output_1_3_0_15_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_19_8_sva <= R_19_6_sva ^ (s_output_1_19_16_41_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_12_8_sva <= R_12_6_sva ^ (s_output_1_19_16_11_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_18_8_sva <= R_18_6_sva ^ (s_output_1_3_0_30_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_13_8_sva <= R_13_6_sva ^ (s_output_1_3_0_45_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_17_8_sva <= R_17_6_sva ^ (s_output_1_3_0_15_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_14_8_sva <= R_14_6_sva ^ (s_output_1_19_16_41_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_16_8_sva <= R_16_6_sva ^ (s_output_1_19_16_56_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[7] ) begin
      R_15_8_sva <= R_15_6_sva ^ (s_output_1_19_16_26_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_31_9_sva <= R_31_7_sva ^ (s_output_1_19_16_12_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_0_9_sva <= R_0_7_sva ^ (s_output_1_3_0_61_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_30_9_sva <= R_30_7_sva ^ (s_output_1_19_16_42_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_1_9_sva <= R_1_7_sva ^ (s_output_1_19_16_27_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_29_9_sva <= R_29_7_sva ^ (s_output_1_3_0_31_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_2_9_sva <= R_2_7_sva ^ (s_output_1_19_16_57_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_28_9_sva <= R_28_7_sva ^ (s_output_1_3_0_46_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_3_9_sva <= R_3_7_sva ^ (s_output_1_3_0_46_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_27_9_sva <= R_27_7_sva ^ (s_output_1_3_0_16_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_4_9_sva <= R_4_7_sva ^ (s_output_1_19_16_42_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_26_9_sva <= R_26_7_sva ^ (s_output_1_19_16_57_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_5_9_sva <= R_5_7_sva ^ (s_output_1_3_0_16_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_25_9_sva <= R_25_7_sva ^ (s_output_1_3_0_61_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_6_9_sva <= R_6_7_sva ^ (s_output_1_19_16_12_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_24_9_sva <= R_24_7_sva ^ (s_output_1_3_0_31_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_7_9_sva <= R_7_7_sva ^ (s_output_1_3_0_31_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_23_9_sva <= R_23_7_sva ^ (s_output_1_19_16_27_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_8_9_sva <= R_8_7_sva ^ (s_output_1_19_16_57_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_22_9_sva <= R_22_7_sva ^ (s_output_1_19_16_12_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_9_9_sva <= R_9_7_sva ^ (s_output_1_19_16_27_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_21_9_sva <= R_21_7_sva ^ (s_output_1_3_0_46_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_10_9_sva <= R_10_7_sva ^ (s_output_1_3_0_61_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_20_9_sva <= R_20_7_sva ^ (s_output_1_3_0_61_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_11_9_sva <= R_11_7_sva ^ (s_output_1_3_0_16_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_19_9_sva <= R_19_7_sva ^ (s_output_1_19_16_42_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_12_9_sva <= R_12_7_sva ^ (s_output_1_19_16_12_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_18_9_sva <= R_18_7_sva ^ (s_output_1_3_0_31_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_13_9_sva <= R_13_7_sva ^ (s_output_1_3_0_46_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_17_9_sva <= R_17_7_sva ^ (s_output_1_3_0_16_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_14_9_sva <= R_14_7_sva ^ (s_output_1_19_16_42_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_16_9_sva <= R_16_7_sva ^ (s_output_1_19_16_57_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[8] ) begin
      R_15_9_sva <= R_15_7_sva ^ (s_output_1_19_16_27_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_31_10_sva <= R_31_8_sva ^ (s_output_1_19_16_13_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_0_10_sva <= R_0_8_sva ^ (s_output_1_3_0_62_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_30_10_sva <= R_30_8_sva ^ (s_output_1_19_16_43_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_1_10_sva <= R_1_8_sva ^ (s_output_1_19_16_28_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_29_10_sva <= R_29_8_sva ^ (s_output_1_3_0_32_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_2_10_sva <= R_2_8_sva ^ (s_output_1_19_16_58_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_28_10_sva <= R_28_8_sva ^ (s_output_1_3_0_47_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_3_10_sva <= R_3_8_sva ^ (s_output_1_3_0_47_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_27_10_sva <= R_27_8_sva ^ (s_output_1_3_0_17_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_4_10_sva <= R_4_8_sva ^ (s_output_1_19_16_43_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_26_10_sva <= R_26_8_sva ^ (s_output_1_19_16_58_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_5_10_sva <= R_5_8_sva ^ (s_output_1_3_0_17_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_25_10_sva <= R_25_8_sva ^ (s_output_1_3_0_62_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_6_10_sva <= R_6_8_sva ^ (s_output_1_19_16_13_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_24_10_sva <= R_24_8_sva ^ (s_output_1_3_0_32_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_7_10_sva <= R_7_8_sva ^ (s_output_1_3_0_32_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_23_10_sva <= R_23_8_sva ^ (s_output_1_19_16_28_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_8_10_sva <= R_8_8_sva ^ (s_output_1_19_16_58_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_22_10_sva <= R_22_8_sva ^ (s_output_1_19_16_13_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_9_10_sva <= R_9_8_sva ^ (s_output_1_19_16_28_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_21_10_sva <= R_21_8_sva ^ (s_output_1_3_0_47_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_10_10_sva <= R_10_8_sva ^ (s_output_1_3_0_62_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_20_10_sva <= R_20_8_sva ^ (s_output_1_3_0_62_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_11_10_sva <= R_11_8_sva ^ (s_output_1_3_0_17_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_19_10_sva <= R_19_8_sva ^ (s_output_1_19_16_43_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_12_10_sva <= R_12_8_sva ^ (s_output_1_19_16_13_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_18_10_sva <= R_18_8_sva ^ (s_output_1_3_0_32_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_13_10_sva <= R_13_8_sva ^ (s_output_1_3_0_47_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_17_10_sva <= R_17_8_sva ^ (s_output_1_3_0_17_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_14_10_sva <= R_14_8_sva ^ (s_output_1_19_16_43_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_16_10_sva <= R_16_8_sva ^ (s_output_1_19_16_58_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[9] ) begin
      R_15_10_sva <= R_15_8_sva ^ (s_output_1_19_16_28_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_31_11_sva <= R_31_9_sva ^ (s_output_1_19_16_14_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_0_11_sva <= R_0_9_sva ^ (s_output_1_3_0_63_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_30_11_sva <= R_30_9_sva ^ (s_output_1_19_16_44_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_1_11_sva <= R_1_9_sva ^ (s_output_1_19_16_29_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_29_11_sva <= R_29_9_sva ^ (s_output_1_3_0_33_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_2_11_sva <= R_2_9_sva ^ (s_output_1_19_16_59_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_28_11_sva <= R_28_9_sva ^ (s_output_1_3_0_48_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_3_11_sva <= R_3_9_sva ^ (s_output_1_3_0_48_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_27_11_sva <= R_27_9_sva ^ (s_output_1_3_0_18_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_4_11_sva <= R_4_9_sva ^ (s_output_1_19_16_44_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_26_11_sva <= R_26_9_sva ^ (s_output_1_19_16_59_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_5_11_sva <= R_5_9_sva ^ (s_output_1_3_0_18_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_25_11_sva <= R_25_9_sva ^ (s_output_1_3_0_63_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_6_11_sva <= R_6_9_sva ^ (s_output_1_19_16_14_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_24_11_sva <= R_24_9_sva ^ (s_output_1_3_0_33_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_7_11_sva <= R_7_9_sva ^ (s_output_1_3_0_33_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_23_11_sva <= R_23_9_sva ^ (s_output_1_19_16_29_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_8_11_sva <= R_8_9_sva ^ (s_output_1_19_16_59_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_22_11_sva <= R_22_9_sva ^ (s_output_1_19_16_14_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_9_11_sva <= R_9_9_sva ^ (s_output_1_19_16_29_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_21_11_sva <= R_21_9_sva ^ (s_output_1_3_0_48_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_10_11_sva <= R_10_9_sva ^ (s_output_1_3_0_63_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_20_11_sva <= R_20_9_sva ^ (s_output_1_3_0_63_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_11_11_sva <= R_11_9_sva ^ (s_output_1_3_0_18_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_19_11_sva <= R_19_9_sva ^ (s_output_1_19_16_44_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_12_11_sva <= R_12_9_sva ^ (s_output_1_19_16_14_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_18_11_sva <= R_18_9_sva ^ (s_output_1_3_0_33_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_13_11_sva <= R_13_9_sva ^ (s_output_1_3_0_48_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_17_11_sva <= R_17_9_sva ^ (s_output_1_3_0_18_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_14_11_sva <= R_14_9_sva ^ (s_output_1_19_16_44_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_16_11_sva <= R_16_9_sva ^ (s_output_1_19_16_59_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[10] ) begin
      R_15_11_sva <= R_15_9_sva ^ (s_output_1_19_16_29_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_31_12_sva <= R_31_10_sva ^ (s_output_1_19_16_15_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_0_12_sva <= R_0_10_sva ^ (s_output_1_3_0_64_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_30_12_sva <= R_30_10_sva ^ (s_output_1_19_16_45_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_1_12_sva <= R_1_10_sva ^ (s_output_1_19_16_30_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_29_12_sva <= R_29_10_sva ^ (s_output_1_3_0_34_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_2_12_sva <= R_2_10_sva ^ (s_output_1_19_16_60_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_28_12_sva <= R_28_10_sva ^ (s_output_1_3_0_49_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_3_12_sva <= R_3_10_sva ^ (s_output_1_3_0_49_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_27_12_sva <= R_27_10_sva ^ (s_output_1_3_0_19_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_4_12_sva <= R_4_10_sva ^ (s_output_1_19_16_45_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_26_12_sva <= R_26_10_sva ^ (s_output_1_19_16_60_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_5_12_sva <= R_5_10_sva ^ (s_output_1_3_0_19_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_25_12_sva <= R_25_10_sva ^ (s_output_1_3_0_64_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_6_12_sva <= R_6_10_sva ^ (s_output_1_19_16_15_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_24_12_sva <= R_24_10_sva ^ (s_output_1_3_0_34_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_7_12_sva <= R_7_10_sva ^ (s_output_1_3_0_34_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_23_12_sva <= R_23_10_sva ^ (s_output_1_19_16_30_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_8_12_sva <= R_8_10_sva ^ (s_output_1_19_16_60_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_22_12_sva <= R_22_10_sva ^ (s_output_1_19_16_15_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_9_12_sva <= R_9_10_sva ^ (s_output_1_19_16_30_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_21_12_sva <= R_21_10_sva ^ (s_output_1_3_0_49_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_10_12_sva <= R_10_10_sva ^ (s_output_1_3_0_64_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_20_12_sva <= R_20_10_sva ^ (s_output_1_3_0_64_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_11_12_sva <= R_11_10_sva ^ (s_output_1_3_0_19_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_19_12_sva <= R_19_10_sva ^ (s_output_1_19_16_45_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_12_12_sva <= R_12_10_sva ^ (s_output_1_19_16_15_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_18_12_sva <= R_18_10_sva ^ (s_output_1_3_0_34_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_13_12_sva <= R_13_10_sva ^ (s_output_1_3_0_49_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_17_12_sva <= R_17_10_sva ^ (s_output_1_3_0_19_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_14_12_sva <= R_14_10_sva ^ (s_output_1_19_16_45_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_16_12_sva <= R_16_10_sva ^ (s_output_1_19_16_60_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[11] ) begin
      R_15_12_sva <= R_15_10_sva ^ (s_output_1_19_16_30_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_31_13_sva <= R_31_11_sva ^ (s_output_1_19_16_16_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_0_13_sva <= R_0_11_sva ^ (s_output_1_3_0_65_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_30_13_sva <= R_30_11_sva ^ (s_output_1_19_16_46_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_1_13_sva <= R_1_11_sva ^ (s_output_1_19_16_31_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_29_13_sva <= R_29_11_sva ^ (s_output_1_3_0_35_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_2_13_sva <= R_2_11_sva ^ (s_output_1_19_16_61_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_28_13_sva <= R_28_11_sva ^ (s_output_1_3_0_50_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_3_13_sva <= R_3_11_sva ^ (s_output_1_3_0_50_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_27_13_sva <= R_27_11_sva ^ (s_output_1_3_0_20_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_4_13_sva <= R_4_11_sva ^ (s_output_1_19_16_46_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_26_13_sva <= R_26_11_sva ^ (s_output_1_19_16_61_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_5_13_sva <= R_5_11_sva ^ (s_output_1_3_0_20_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_25_13_sva <= R_25_11_sva ^ (s_output_1_3_0_65_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_6_13_sva <= R_6_11_sva ^ (s_output_1_19_16_16_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_24_13_sva <= R_24_11_sva ^ (s_output_1_3_0_35_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_7_13_sva <= R_7_11_sva ^ (s_output_1_3_0_35_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_23_13_sva <= R_23_11_sva ^ (s_output_1_19_16_31_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_8_13_sva <= R_8_11_sva ^ (s_output_1_19_16_61_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_22_13_sva <= R_22_11_sva ^ (s_output_1_19_16_16_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_9_13_sva <= R_9_11_sva ^ (s_output_1_19_16_31_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_21_13_sva <= R_21_11_sva ^ (s_output_1_3_0_50_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_10_13_sva <= R_10_11_sva ^ (s_output_1_3_0_65_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_20_13_sva <= R_20_11_sva ^ (s_output_1_3_0_65_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_11_13_sva <= R_11_11_sva ^ (s_output_1_3_0_20_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_19_13_sva <= R_19_11_sva ^ (s_output_1_19_16_46_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_12_13_sva <= R_12_11_sva ^ (s_output_1_19_16_16_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_18_13_sva <= R_18_11_sva ^ (s_output_1_3_0_35_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_13_13_sva <= R_13_11_sva ^ (s_output_1_3_0_50_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_17_13_sva <= R_17_11_sva ^ (s_output_1_3_0_20_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_14_13_sva <= R_14_11_sva ^ (s_output_1_19_16_46_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_16_13_sva <= R_16_11_sva ^ (s_output_1_19_16_61_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[12] ) begin
      R_15_13_sva <= R_15_11_sva ^ (s_output_1_19_16_31_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_7_14_sva <= R_7_12_sva ^ (s_output_1_3_0_36_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_24_14_sva <= R_24_12_sva ^ (s_output_1_3_0_36_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_15_14_sva <= R_15_12_sva ^ (s_output_1_19_16_32_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_16_14_sva <= R_16_12_sva ^ (s_output_1_19_16_62_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_23_14_sva <= R_23_12_sva ^ (s_output_1_19_16_32_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_8_14_sva <= R_8_12_sva ^ (s_output_1_19_16_62_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_31_14_sva <= R_31_12_sva ^ (s_output_1_19_16_17_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_0_14_sva <= R_0_12_sva ^ (s_output_1_3_0_66_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_6_14_sva <= R_6_12_sva ^ (s_output_1_19_16_17_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_25_14_sva <= R_25_12_sva ^ (s_output_1_3_0_66_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_14_14_sva <= R_14_12_sva ^ (s_output_1_19_16_47_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_17_14_sva <= R_17_12_sva ^ (s_output_1_3_0_21_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_22_14_sva <= R_22_12_sva ^ (s_output_1_19_16_17_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_9_14_sva <= R_9_12_sva ^ (s_output_1_19_16_32_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_30_14_sva <= R_30_12_sva ^ (s_output_1_19_16_47_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_1_14_sva <= R_1_12_sva ^ (s_output_1_19_16_32_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_5_14_sva <= R_5_12_sva ^ (s_output_1_3_0_21_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_26_14_sva <= R_26_12_sva ^ (s_output_1_19_16_62_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_13_14_sva <= R_13_12_sva ^ (s_output_1_3_0_51_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_18_14_sva <= R_18_12_sva ^ (s_output_1_3_0_36_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_21_14_sva <= R_21_12_sva ^ (s_output_1_3_0_51_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_10_14_sva <= R_10_12_sva ^ (s_output_1_3_0_66_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_29_14_sva <= R_29_12_sva ^ (s_output_1_3_0_36_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_2_14_sva <= R_2_12_sva ^ (s_output_1_19_16_62_sva_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_4_14_sva <= R_4_12_sva ^ (s_output_1_19_16_47_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_27_14_sva <= R_27_12_sva ^ (s_output_1_3_0_21_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_12_14_sva <= R_12_12_sva ^ (s_output_1_19_16_17_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_19_14_sva <= R_19_12_sva ^ (s_output_1_19_16_47_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_20_14_sva <= R_20_12_sva ^ (s_output_1_3_0_66_sva_1[2]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_11_14_sva <= R_11_12_sva ^ (s_output_1_3_0_21_sva_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_28_14_sva <= R_28_12_sva ^ (s_output_1_3_0_51_sva_1[3]);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[13] ) begin
      R_3_14_sva <= R_3_12_sva ^ (s_output_1_3_0_51_sva_1[2]);
    end
  end
  assign loop_DES_rounds_1_xor_32_nl = (input_sva[6]) ^ (s_output_1_19_16_4_sva[0]);
  assign loop_DES_rounds_2_xor_32_nl = (input_sva[7]) ^ (s_output_1_19_16_5_sva[0]);
  assign loop_DES_rounds_1_xor_31_nl = (input_sva[56]) ^ (s_output_1_3_0_53_sva[3]);
  assign loop_DES_rounds_2_xor_31_nl = (input_sva[57]) ^ (s_output_1_3_0_54_sva[3]);
  assign loop_DES_rounds_1_xor_30_nl = (input_sva[14]) ^ (s_output_1_19_16_34_sva[1]);
  assign loop_DES_rounds_2_xor_30_nl = (input_sva[15]) ^ (s_output_1_19_16_35_sva[1]);
  assign loop_DES_rounds_1_xor_29_nl = (input_sva[48]) ^ (s_output_1_19_16_19_sva[0]);
  assign loop_DES_rounds_2_xor_29_nl = (input_sva[49]) ^ (s_output_1_19_16_20_sva[0]);
  assign loop_DES_rounds_1_xor_28_nl = (input_sva[22]) ^ (s_output_1_3_0_23_sva[0]);
  assign loop_DES_rounds_2_xor_28_nl = (input_sva[23]) ^ (s_output_1_3_0_24_sva[0]);
  assign loop_DES_rounds_1_xor_27_nl = (input_sva[40]) ^ (s_output_1_19_16_49_sva[1]);
  assign loop_DES_rounds_2_xor_27_nl = (input_sva[41]) ^ (s_output_1_19_16_50_sva[1]);
  assign loop_DES_rounds_1_xor_26_nl = (input_sva[30]) ^ (s_output_1_3_0_38_sva[3]);
  assign loop_DES_rounds_2_xor_26_nl = (input_sva[31]) ^ (s_output_1_3_0_39_sva[3]);
  assign loop_DES_rounds_1_xor_25_nl = (input_sva[32]) ^ (s_output_1_3_0_38_sva[2]);
  assign loop_DES_rounds_2_xor_25_nl = (input_sva[33]) ^ (s_output_1_3_0_39_sva[2]);
  assign loop_DES_rounds_1_xor_24_nl = (input_sva[38]) ^ (s_output_1_3_0_8_sva[3]);
  assign loop_DES_rounds_2_xor_24_nl = (input_sva[39]) ^ (s_output_1_3_0_9_sva[3]);
  assign loop_DES_rounds_1_xor_23_nl = (input_sva[24]) ^ (s_output_1_19_16_34_sva[2]);
  assign loop_DES_rounds_2_xor_23_nl = (input_sva[25]) ^ (s_output_1_19_16_35_sva[2]);
  assign loop_DES_rounds_1_xor_22_nl = (input_sva[46]) ^ (s_output_1_19_16_49_sva[0]);
  assign loop_DES_rounds_2_xor_22_nl = (input_sva[47]) ^ (s_output_1_19_16_50_sva[0]);
  assign loop_DES_rounds_1_xor_21_nl = (input_sva[16]) ^ (s_output_1_3_0_8_sva[2]);
  assign loop_DES_rounds_2_xor_21_nl = (input_sva[17]) ^ (s_output_1_3_0_9_sva[2]);
  assign loop_DES_rounds_1_xor_20_nl = (input_sva[54]) ^ (s_output_1_3_0_53_sva[0]);
  assign loop_DES_rounds_2_xor_20_nl = (input_sva[55]) ^ (s_output_1_3_0_54_sva[0]);
  assign loop_DES_rounds_1_xor_19_nl = (input_sva[8]) ^ (s_output_1_19_16_4_sva[3]);
  assign loop_DES_rounds_2_xor_19_nl = (input_sva[9]) ^ (s_output_1_19_16_5_sva[3]);
  assign loop_DES_rounds_1_xor_18_nl = (input_sva[62]) ^ (s_output_1_3_0_23_sva[3]);
  assign loop_DES_rounds_2_xor_18_nl = (input_sva[63]) ^ (s_output_1_3_0_24_sva[3]);
  assign loop_DES_rounds_1_xor_17_nl = (input_sva[0]) ^ (s_output_1_3_0_23_sva[1]);
  assign loop_DES_rounds_2_xor_17_nl = (input_sva[1]) ^ (s_output_1_3_0_24_sva[1]);
  assign loop_DES_rounds_1_xor_16_nl = (input_sva[4]) ^ (s_output_1_19_16_19_sva[3]);
  assign loop_DES_rounds_2_xor_16_nl = (input_sva[5]) ^ (s_output_1_19_16_20_sva[3]);
  assign loop_DES_rounds_1_xor_15_nl = (input_sva[58]) ^ (s_output_1_19_16_49_sva[3]);
  assign loop_DES_rounds_2_xor_15_nl = (input_sva[59]) ^ (s_output_1_19_16_50_sva[3]);
  assign loop_DES_rounds_1_xor_14_nl = (input_sva[12]) ^ (s_output_1_19_16_4_sva[1]);
  assign loop_DES_rounds_2_xor_14_nl = (input_sva[13]) ^ (s_output_1_19_16_5_sva[1]);
  assign loop_DES_rounds_1_xor_13_nl = (input_sva[50]) ^ (s_output_1_19_16_19_sva[1]);
  assign loop_DES_rounds_2_xor_13_nl = (input_sva[51]) ^ (s_output_1_19_16_20_sva[1]);
  assign loop_DES_rounds_1_xor_12_nl = (input_sva[20]) ^ (s_output_1_3_0_38_sva[1]);
  assign loop_DES_rounds_2_xor_12_nl = (input_sva[21]) ^ (s_output_1_3_0_39_sva[1]);
  assign loop_DES_rounds_1_xor_11_nl = (input_sva[42]) ^ (s_output_1_3_0_53_sva[1]);
  assign loop_DES_rounds_2_xor_11_nl = (input_sva[43]) ^ (s_output_1_3_0_54_sva[1]);
  assign loop_DES_rounds_1_xor_10_nl = (input_sva[28]) ^ (s_output_1_3_0_53_sva[2]);
  assign loop_DES_rounds_2_xor_10_nl = (input_sva[29]) ^ (s_output_1_3_0_54_sva[2]);
  assign loop_DES_rounds_1_xor_9_nl = (input_sva[34]) ^ (s_output_1_3_0_8_sva[0]);
  assign loop_DES_rounds_2_xor_9_nl = (input_sva[35]) ^ (s_output_1_3_0_9_sva[0]);
  assign loop_DES_rounds_1_xor_8_nl = (input_sva[36]) ^ (s_output_1_19_16_34_sva[3]);
  assign loop_DES_rounds_2_xor_8_nl = (input_sva[37]) ^ (s_output_1_19_16_35_sva[3]);
  assign loop_DES_rounds_1_xor_7_nl = (input_sva[26]) ^ (s_output_1_19_16_4_sva[2]);
  assign loop_DES_rounds_2_xor_7_nl = (input_sva[27]) ^ (s_output_1_19_16_5_sva[2]);
  assign loop_DES_rounds_1_xor_6_nl = (input_sva[44]) ^ (s_output_1_3_0_23_sva[2]);
  assign loop_DES_rounds_2_xor_6_nl = (input_sva[45]) ^ (s_output_1_3_0_24_sva[2]);
  assign loop_DES_rounds_1_xor_5_nl = (input_sva[18]) ^ (s_output_1_3_0_38_sva[0]);
  assign loop_DES_rounds_2_xor_5_nl = (input_sva[19]) ^ (s_output_1_3_0_39_sva[0]);
  assign loop_DES_rounds_1_xor_4_nl = (input_sva[52]) ^ (s_output_1_3_0_8_sva[1]);
  assign loop_DES_rounds_2_xor_4_nl = (input_sva[53]) ^ (s_output_1_3_0_9_sva[1]);
  assign loop_DES_rounds_1_xor_3_nl = (input_sva[10]) ^ (s_output_1_19_16_34_sva[0]);
  assign loop_DES_rounds_2_xor_3_nl = (input_sva[11]) ^ (s_output_1_19_16_35_sva[0]);
  assign loop_DES_rounds_1_xor_2_nl = (input_sva[60]) ^ (s_output_1_19_16_49_sva[2]);
  assign loop_DES_rounds_2_xor_2_nl = (input_sva[61]) ^ (s_output_1_19_16_50_sva[2]);
  assign loop_DES_rounds_1_xor_1_nl = (input_sva[2]) ^ (s_output_1_19_16_19_sva[2]);
  assign loop_DES_rounds_2_xor_1_nl = (input_sva[3]) ^ (s_output_1_19_16_20_sva[2]);

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    des_check
// ------------------------------------------------------------------


module des_check (
  clk, rst, input_rsc_dat, input_rsc_triosy_lz, key_rsc_dat, key_rsc_triosy_lz, return_rsc_dat,
      return_rsc_triosy_lz
);
  input clk;
  input rst;
  input [63:0] input_rsc_dat;
  output input_rsc_triosy_lz;
  input [63:0] key_rsc_dat;
  output key_rsc_triosy_lz;
  output [63:0] return_rsc_dat;
  output return_rsc_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  des_check_core des_check_core_inst (
      .clk(clk),
      .rst(rst),
      .input_rsc_dat(input_rsc_dat),
      .input_rsc_triosy_lz(input_rsc_triosy_lz),
      .key_rsc_dat(key_rsc_dat),
      .key_rsc_triosy_lz(key_rsc_triosy_lz),
      .return_rsc_dat(return_rsc_dat),
      .return_rsc_triosy_lz(return_rsc_triosy_lz)
    );
endmodule



