
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ../td_ccore_solutions/ROM_1i6_1o4_cfafff97e973ca9580e646fecdc2f814b3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Mon Mar  1 00:26:13 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i6_1o4_cfafff97e973ca9580e646fecdc2f814b3
// ------------------------------------------------------------------


module ROM_1i6_1o4_cfafff97e973ca9580e646fecdc2f814b3 (
  I_1, O_1
);
  input [5:0] I_1;
  output [3:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_4_64_2(4'b1111, 4'b0001, 4'b1000, 4'b1110, 4'b0110, 4'b1011,
      4'b0011, 4'b0100, 4'b1001, 4'b0111, 4'b0010, 4'b1101, 4'b1100, 4'b0000, 4'b0101,
      4'b1010, 4'b0011, 4'b1101, 4'b0100, 4'b0111, 4'b1111, 4'b0010, 4'b1000, 4'b1110,
      4'b1100, 4'b0000, 4'b0001, 4'b1010, 4'b0110, 4'b1001, 4'b1011, 4'b0101, 4'b0000,
      4'b1110, 4'b0111, 4'b1011, 4'b1010, 4'b0100, 4'b1101, 4'b0001, 4'b0101, 4'b1000,
      4'b1100, 4'b0110, 4'b1001, 4'b0011, 4'b0010, 4'b1111, 4'b1101, 4'b1000, 4'b1010,
      4'b0001, 4'b0011, 4'b1111, 4'b0100, 4'b0010, 4'b1011, 4'b0110, 4'b0111, 4'b1100,
      4'b0000, 4'b0101, 4'b1110, 4'b1001, I_1);

  function automatic [3:0] MUX_v_4_64_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [3:0] input_8;
    input [3:0] input_9;
    input [3:0] input_10;
    input [3:0] input_11;
    input [3:0] input_12;
    input [3:0] input_13;
    input [3:0] input_14;
    input [3:0] input_15;
    input [3:0] input_16;
    input [3:0] input_17;
    input [3:0] input_18;
    input [3:0] input_19;
    input [3:0] input_20;
    input [3:0] input_21;
    input [3:0] input_22;
    input [3:0] input_23;
    input [3:0] input_24;
    input [3:0] input_25;
    input [3:0] input_26;
    input [3:0] input_27;
    input [3:0] input_28;
    input [3:0] input_29;
    input [3:0] input_30;
    input [3:0] input_31;
    input [3:0] input_32;
    input [3:0] input_33;
    input [3:0] input_34;
    input [3:0] input_35;
    input [3:0] input_36;
    input [3:0] input_37;
    input [3:0] input_38;
    input [3:0] input_39;
    input [3:0] input_40;
    input [3:0] input_41;
    input [3:0] input_42;
    input [3:0] input_43;
    input [3:0] input_44;
    input [3:0] input_45;
    input [3:0] input_46;
    input [3:0] input_47;
    input [3:0] input_48;
    input [3:0] input_49;
    input [3:0] input_50;
    input [3:0] input_51;
    input [3:0] input_52;
    input [3:0] input_53;
    input [3:0] input_54;
    input [3:0] input_55;
    input [3:0] input_56;
    input [3:0] input_57;
    input [3:0] input_58;
    input [3:0] input_59;
    input [3:0] input_60;
    input [3:0] input_61;
    input [3:0] input_62;
    input [3:0] input_63;
    input [5:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_4_64_2 = result;
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i6_1o4_d0e242163cbb0b2ce9c4399bc1cb50f5b3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Mon Mar  1 00:26:47 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i6_1o4_d0e242163cbb0b2ce9c4399bc1cb50f5b3
// ------------------------------------------------------------------


module ROM_1i6_1o4_d0e242163cbb0b2ce9c4399bc1cb50f5b3 (
  I_1, O_1
);
  input [5:0] I_1;
  output [3:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_4_64_2(4'b0111, 4'b1101, 4'b1110, 4'b0011, 4'b0000, 4'b0110,
      4'b1001, 4'b1010, 4'b0001, 4'b0010, 4'b1000, 4'b0101, 4'b1011, 4'b1100, 4'b0100,
      4'b1111, 4'b1101, 4'b1000, 4'b1011, 4'b0101, 4'b0110, 4'b1111, 4'b0000, 4'b0011,
      4'b0100, 4'b0111, 4'b0010, 4'b1100, 4'b0001, 4'b1010, 4'b1110, 4'b1001, 4'b1010,
      4'b0110, 4'b1001, 4'b0000, 4'b1100, 4'b1011, 4'b0111, 4'b1101, 4'b1111, 4'b0001,
      4'b0011, 4'b1110, 4'b0101, 4'b0010, 4'b1000, 4'b0100, 4'b0011, 4'b1111, 4'b0000,
      4'b0110, 4'b1010, 4'b0001, 4'b1101, 4'b1000, 4'b1001, 4'b0100, 4'b0101, 4'b1011,
      4'b1100, 4'b0111, 4'b0010, 4'b1110, I_1);

  function automatic [3:0] MUX_v_4_64_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [3:0] input_8;
    input [3:0] input_9;
    input [3:0] input_10;
    input [3:0] input_11;
    input [3:0] input_12;
    input [3:0] input_13;
    input [3:0] input_14;
    input [3:0] input_15;
    input [3:0] input_16;
    input [3:0] input_17;
    input [3:0] input_18;
    input [3:0] input_19;
    input [3:0] input_20;
    input [3:0] input_21;
    input [3:0] input_22;
    input [3:0] input_23;
    input [3:0] input_24;
    input [3:0] input_25;
    input [3:0] input_26;
    input [3:0] input_27;
    input [3:0] input_28;
    input [3:0] input_29;
    input [3:0] input_30;
    input [3:0] input_31;
    input [3:0] input_32;
    input [3:0] input_33;
    input [3:0] input_34;
    input [3:0] input_35;
    input [3:0] input_36;
    input [3:0] input_37;
    input [3:0] input_38;
    input [3:0] input_39;
    input [3:0] input_40;
    input [3:0] input_41;
    input [3:0] input_42;
    input [3:0] input_43;
    input [3:0] input_44;
    input [3:0] input_45;
    input [3:0] input_46;
    input [3:0] input_47;
    input [3:0] input_48;
    input [3:0] input_49;
    input [3:0] input_50;
    input [3:0] input_51;
    input [3:0] input_52;
    input [3:0] input_53;
    input [3:0] input_54;
    input [3:0] input_55;
    input [3:0] input_56;
    input [3:0] input_57;
    input [3:0] input_58;
    input [3:0] input_59;
    input [3:0] input_60;
    input [3:0] input_61;
    input [3:0] input_62;
    input [3:0] input_63;
    input [5:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_4_64_2 = result;
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i6_1o4_752c7ca65a598ada4acee0cd63d199c3b3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Mon Mar  1 00:26:38 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i6_1o4_752c7ca65a598ada4acee0cd63d199c3b3
// ------------------------------------------------------------------


module ROM_1i6_1o4_752c7ca65a598ada4acee0cd63d199c3b3 (
  I_1, O_1
);
  input [5:0] I_1;
  output [3:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_4_64_2(4'b0100, 4'b1011, 4'b0010, 4'b1110, 4'b1111, 4'b0000,
      4'b1000, 4'b1101, 4'b0011, 4'b1100, 4'b1001, 4'b0111, 4'b0101, 4'b1010, 4'b0110,
      4'b0001, 4'b1101, 4'b0000, 4'b1011, 4'b0111, 4'b0100, 4'b1001, 4'b0001, 4'b1010,
      4'b1110, 4'b0011, 4'b0101, 4'b1100, 4'b0010, 4'b1111, 4'b1000, 4'b0110, 4'b0001,
      4'b0100, 4'b1011, 4'b1101, 4'b1100, 4'b0011, 4'b0111, 4'b1110, 4'b1010, 4'b1111,
      4'b0110, 4'b1000, 4'b0000, 4'b0101, 4'b1001, 4'b0010, 4'b0110, 4'b1011, 4'b1101,
      4'b1000, 4'b0001, 4'b0100, 4'b1010, 4'b0111, 4'b1001, 4'b0101, 4'b0000, 4'b1111,
      4'b1110, 4'b0010, 4'b0011, 4'b1100, I_1);

  function automatic [3:0] MUX_v_4_64_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [3:0] input_8;
    input [3:0] input_9;
    input [3:0] input_10;
    input [3:0] input_11;
    input [3:0] input_12;
    input [3:0] input_13;
    input [3:0] input_14;
    input [3:0] input_15;
    input [3:0] input_16;
    input [3:0] input_17;
    input [3:0] input_18;
    input [3:0] input_19;
    input [3:0] input_20;
    input [3:0] input_21;
    input [3:0] input_22;
    input [3:0] input_23;
    input [3:0] input_24;
    input [3:0] input_25;
    input [3:0] input_26;
    input [3:0] input_27;
    input [3:0] input_28;
    input [3:0] input_29;
    input [3:0] input_30;
    input [3:0] input_31;
    input [3:0] input_32;
    input [3:0] input_33;
    input [3:0] input_34;
    input [3:0] input_35;
    input [3:0] input_36;
    input [3:0] input_37;
    input [3:0] input_38;
    input [3:0] input_39;
    input [3:0] input_40;
    input [3:0] input_41;
    input [3:0] input_42;
    input [3:0] input_43;
    input [3:0] input_44;
    input [3:0] input_45;
    input [3:0] input_46;
    input [3:0] input_47;
    input [3:0] input_48;
    input [3:0] input_49;
    input [3:0] input_50;
    input [3:0] input_51;
    input [3:0] input_52;
    input [3:0] input_53;
    input [3:0] input_54;
    input [3:0] input_55;
    input [3:0] input_56;
    input [3:0] input_57;
    input [3:0] input_58;
    input [3:0] input_59;
    input [3:0] input_60;
    input [3:0] input_61;
    input [3:0] input_62;
    input [3:0] input_63;
    input [5:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_4_64_2 = result;
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i6_1o4_ef717c7c87dc90ac6f7b34d533fe115fb3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Mon Mar  1 00:26:05 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i6_1o4_ef717c7c87dc90ac6f7b34d533fe115fb3
// ------------------------------------------------------------------


module ROM_1i6_1o4_ef717c7c87dc90ac6f7b34d533fe115fb3 (
  I_1, O_1
);
  input [5:0] I_1;
  output [3:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_4_64_2(4'b0010, 4'b1100, 4'b0100, 4'b0001, 4'b0111, 4'b1010,
      4'b1011, 4'b0110, 4'b1000, 4'b0101, 4'b0011, 4'b1111, 4'b1101, 4'b0000, 4'b1110,
      4'b1001, 4'b1110, 4'b1011, 4'b0010, 4'b1100, 4'b0100, 4'b0111, 4'b1101, 4'b0001,
      4'b0101, 4'b0000, 4'b1111, 4'b1010, 4'b0011, 4'b1001, 4'b1000, 4'b0110, 4'b0100,
      4'b0010, 4'b0001, 4'b1011, 4'b1010, 4'b1101, 4'b0111, 4'b1000, 4'b1111, 4'b1001,
      4'b1100, 4'b0101, 4'b0110, 4'b0011, 4'b0000, 4'b1110, 4'b1011, 4'b1000, 4'b1100,
      4'b0111, 4'b0001, 4'b1110, 4'b0010, 4'b1101, 4'b0110, 4'b1111, 4'b0000, 4'b1001,
      4'b1010, 4'b0100, 4'b0101, 4'b0011, I_1);

  function automatic [3:0] MUX_v_4_64_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [3:0] input_8;
    input [3:0] input_9;
    input [3:0] input_10;
    input [3:0] input_11;
    input [3:0] input_12;
    input [3:0] input_13;
    input [3:0] input_14;
    input [3:0] input_15;
    input [3:0] input_16;
    input [3:0] input_17;
    input [3:0] input_18;
    input [3:0] input_19;
    input [3:0] input_20;
    input [3:0] input_21;
    input [3:0] input_22;
    input [3:0] input_23;
    input [3:0] input_24;
    input [3:0] input_25;
    input [3:0] input_26;
    input [3:0] input_27;
    input [3:0] input_28;
    input [3:0] input_29;
    input [3:0] input_30;
    input [3:0] input_31;
    input [3:0] input_32;
    input [3:0] input_33;
    input [3:0] input_34;
    input [3:0] input_35;
    input [3:0] input_36;
    input [3:0] input_37;
    input [3:0] input_38;
    input [3:0] input_39;
    input [3:0] input_40;
    input [3:0] input_41;
    input [3:0] input_42;
    input [3:0] input_43;
    input [3:0] input_44;
    input [3:0] input_45;
    input [3:0] input_46;
    input [3:0] input_47;
    input [3:0] input_48;
    input [3:0] input_49;
    input [3:0] input_50;
    input [3:0] input_51;
    input [3:0] input_52;
    input [3:0] input_53;
    input [3:0] input_54;
    input [3:0] input_55;
    input [3:0] input_56;
    input [3:0] input_57;
    input [3:0] input_58;
    input [3:0] input_59;
    input [3:0] input_60;
    input [3:0] input_61;
    input [3:0] input_62;
    input [3:0] input_63;
    input [5:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_4_64_2 = result;
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i6_1o4_3c5c29b75c561d2b741f22e5a3a569dbb3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Mon Mar  1 00:26:30 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i6_1o4_3c5c29b75c561d2b741f22e5a3a569dbb3
// ------------------------------------------------------------------


module ROM_1i6_1o4_3c5c29b75c561d2b741f22e5a3a569dbb3 (
  I_1, O_1
);
  input [5:0] I_1;
  output [3:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_4_64_2(4'b1010, 4'b0000, 4'b1001, 4'b1110, 4'b0110, 4'b0011,
      4'b1111, 4'b0101, 4'b0001, 4'b1101, 4'b1100, 4'b0111, 4'b1011, 4'b0100, 4'b0010,
      4'b1000, 4'b1101, 4'b0111, 4'b0000, 4'b1001, 4'b0011, 4'b0100, 4'b0110, 4'b1010,
      4'b0010, 4'b1000, 4'b0101, 4'b1110, 4'b1100, 4'b1011, 4'b1111, 4'b0001, 4'b1101,
      4'b0110, 4'b0100, 4'b1001, 4'b1000, 4'b1111, 4'b0011, 4'b0000, 4'b1011, 4'b0001,
      4'b0010, 4'b1100, 4'b0101, 4'b1010, 4'b1110, 4'b0111, 4'b0001, 4'b1010, 4'b1101,
      4'b0000, 4'b0110, 4'b1001, 4'b1000, 4'b0111, 4'b0100, 4'b1111, 4'b1110, 4'b0011,
      4'b1011, 4'b0101, 4'b0010, 4'b1100, I_1);

  function automatic [3:0] MUX_v_4_64_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [3:0] input_8;
    input [3:0] input_9;
    input [3:0] input_10;
    input [3:0] input_11;
    input [3:0] input_12;
    input [3:0] input_13;
    input [3:0] input_14;
    input [3:0] input_15;
    input [3:0] input_16;
    input [3:0] input_17;
    input [3:0] input_18;
    input [3:0] input_19;
    input [3:0] input_20;
    input [3:0] input_21;
    input [3:0] input_22;
    input [3:0] input_23;
    input [3:0] input_24;
    input [3:0] input_25;
    input [3:0] input_26;
    input [3:0] input_27;
    input [3:0] input_28;
    input [3:0] input_29;
    input [3:0] input_30;
    input [3:0] input_31;
    input [3:0] input_32;
    input [3:0] input_33;
    input [3:0] input_34;
    input [3:0] input_35;
    input [3:0] input_36;
    input [3:0] input_37;
    input [3:0] input_38;
    input [3:0] input_39;
    input [3:0] input_40;
    input [3:0] input_41;
    input [3:0] input_42;
    input [3:0] input_43;
    input [3:0] input_44;
    input [3:0] input_45;
    input [3:0] input_46;
    input [3:0] input_47;
    input [3:0] input_48;
    input [3:0] input_49;
    input [3:0] input_50;
    input [3:0] input_51;
    input [3:0] input_52;
    input [3:0] input_53;
    input [3:0] input_54;
    input [3:0] input_55;
    input [3:0] input_56;
    input [3:0] input_57;
    input [3:0] input_58;
    input [3:0] input_59;
    input [3:0] input_60;
    input [3:0] input_61;
    input [3:0] input_62;
    input [3:0] input_63;
    input [5:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_4_64_2 = result;
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i6_1o4_ef4da7ff735c86ba85f23e51741d972cb3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Mon Mar  1 00:26:55 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i6_1o4_ef4da7ff735c86ba85f23e51741d972cb3
// ------------------------------------------------------------------


module ROM_1i6_1o4_ef4da7ff735c86ba85f23e51741d972cb3 (
  I_1, O_1
);
  input [5:0] I_1;
  output [3:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_4_64_2(4'b1101, 4'b0010, 4'b1000, 4'b0100, 4'b0110, 4'b1111,
      4'b1011, 4'b0001, 4'b1010, 4'b1001, 4'b0011, 4'b1110, 4'b0101, 4'b0000, 4'b1100,
      4'b0111, 4'b0001, 4'b1111, 4'b1101, 4'b1000, 4'b1010, 4'b0011, 4'b0111, 4'b0100,
      4'b1100, 4'b0101, 4'b0110, 4'b1011, 4'b0000, 4'b1110, 4'b1001, 4'b0010, 4'b0111,
      4'b1011, 4'b0100, 4'b0001, 4'b1001, 4'b1100, 4'b1110, 4'b0010, 4'b0000, 4'b0110,
      4'b1010, 4'b1101, 4'b1111, 4'b0011, 4'b0101, 4'b1000, 4'b0010, 4'b0001, 4'b1110,
      4'b0111, 4'b0100, 4'b1010, 4'b1000, 4'b1101, 4'b1111, 4'b1100, 4'b1001, 4'b0000,
      4'b0011, 4'b0101, 4'b0110, 4'b1011, I_1);

  function automatic [3:0] MUX_v_4_64_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [3:0] input_8;
    input [3:0] input_9;
    input [3:0] input_10;
    input [3:0] input_11;
    input [3:0] input_12;
    input [3:0] input_13;
    input [3:0] input_14;
    input [3:0] input_15;
    input [3:0] input_16;
    input [3:0] input_17;
    input [3:0] input_18;
    input [3:0] input_19;
    input [3:0] input_20;
    input [3:0] input_21;
    input [3:0] input_22;
    input [3:0] input_23;
    input [3:0] input_24;
    input [3:0] input_25;
    input [3:0] input_26;
    input [3:0] input_27;
    input [3:0] input_28;
    input [3:0] input_29;
    input [3:0] input_30;
    input [3:0] input_31;
    input [3:0] input_32;
    input [3:0] input_33;
    input [3:0] input_34;
    input [3:0] input_35;
    input [3:0] input_36;
    input [3:0] input_37;
    input [3:0] input_38;
    input [3:0] input_39;
    input [3:0] input_40;
    input [3:0] input_41;
    input [3:0] input_42;
    input [3:0] input_43;
    input [3:0] input_44;
    input [3:0] input_45;
    input [3:0] input_46;
    input [3:0] input_47;
    input [3:0] input_48;
    input [3:0] input_49;
    input [3:0] input_50;
    input [3:0] input_51;
    input [3:0] input_52;
    input [3:0] input_53;
    input [3:0] input_54;
    input [3:0] input_55;
    input [3:0] input_56;
    input [3:0] input_57;
    input [3:0] input_58;
    input [3:0] input_59;
    input [3:0] input_60;
    input [3:0] input_61;
    input [3:0] input_62;
    input [3:0] input_63;
    input [5:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_4_64_2 = result;
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i6_1o4_51ba7157b272cd3b87451219caf38e7cb3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Mon Mar  1 00:26:22 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i6_1o4_51ba7157b272cd3b87451219caf38e7cb3
// ------------------------------------------------------------------


module ROM_1i6_1o4_51ba7157b272cd3b87451219caf38e7cb3 (
  I_1, O_1
);
  input [5:0] I_1;
  output [3:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_4_64_2(4'b1100, 4'b0001, 4'b1010, 4'b1111, 4'b1001, 4'b0010,
      4'b0110, 4'b1000, 4'b0000, 4'b1101, 4'b0011, 4'b0100, 4'b1110, 4'b0111, 4'b0101,
      4'b1011, 4'b1010, 4'b1111, 4'b0100, 4'b0010, 4'b0111, 4'b1100, 4'b1001, 4'b0101,
      4'b0110, 4'b0001, 4'b1101, 4'b1110, 4'b0000, 4'b1011, 4'b0011, 4'b1000, 4'b1001,
      4'b1110, 4'b1111, 4'b0101, 4'b0010, 4'b1000, 4'b1100, 4'b0011, 4'b0111, 4'b0000,
      4'b0100, 4'b1010, 4'b0001, 4'b1101, 4'b1011, 4'b0110, 4'b0100, 4'b0011, 4'b0010,
      4'b1100, 4'b1001, 4'b0101, 4'b1111, 4'b1010, 4'b1011, 4'b1110, 4'b0001, 4'b0111,
      4'b0110, 4'b0000, 4'b1000, 4'b1101, I_1);

  function automatic [3:0] MUX_v_4_64_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [3:0] input_8;
    input [3:0] input_9;
    input [3:0] input_10;
    input [3:0] input_11;
    input [3:0] input_12;
    input [3:0] input_13;
    input [3:0] input_14;
    input [3:0] input_15;
    input [3:0] input_16;
    input [3:0] input_17;
    input [3:0] input_18;
    input [3:0] input_19;
    input [3:0] input_20;
    input [3:0] input_21;
    input [3:0] input_22;
    input [3:0] input_23;
    input [3:0] input_24;
    input [3:0] input_25;
    input [3:0] input_26;
    input [3:0] input_27;
    input [3:0] input_28;
    input [3:0] input_29;
    input [3:0] input_30;
    input [3:0] input_31;
    input [3:0] input_32;
    input [3:0] input_33;
    input [3:0] input_34;
    input [3:0] input_35;
    input [3:0] input_36;
    input [3:0] input_37;
    input [3:0] input_38;
    input [3:0] input_39;
    input [3:0] input_40;
    input [3:0] input_41;
    input [3:0] input_42;
    input [3:0] input_43;
    input [3:0] input_44;
    input [3:0] input_45;
    input [3:0] input_46;
    input [3:0] input_47;
    input [3:0] input_48;
    input [3:0] input_49;
    input [3:0] input_50;
    input [3:0] input_51;
    input [3:0] input_52;
    input [3:0] input_53;
    input [3:0] input_54;
    input [3:0] input_55;
    input [3:0] input_56;
    input [3:0] input_57;
    input [3:0] input_58;
    input [3:0] input_59;
    input [3:0] input_60;
    input [3:0] input_61;
    input [3:0] input_62;
    input [3:0] input_63;
    input [5:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_4_64_2 = result;
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i6_1o4_8f60b2fc4a3ee4cef30040071bc0219cb3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Mon Mar  1 00:25:55 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i6_1o4_8f60b2fc4a3ee4cef30040071bc0219cb3
// ------------------------------------------------------------------


module ROM_1i6_1o4_8f60b2fc4a3ee4cef30040071bc0219cb3 (
  I_1, O_1
);
  input [5:0] I_1;
  output [3:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_4_64_2(4'b1110, 4'b0100, 4'b1101, 4'b0001, 4'b0010, 4'b1111,
      4'b1011, 4'b1000, 4'b0011, 4'b1010, 4'b0110, 4'b1100, 4'b0101, 4'b1001, 4'b0000,
      4'b0111, 4'b0000, 4'b1111, 4'b0111, 4'b0100, 4'b1110, 4'b0010, 4'b1101, 4'b0001,
      4'b1010, 4'b0110, 4'b1100, 4'b1011, 4'b1001, 4'b0101, 4'b0011, 4'b1000, 4'b0100,
      4'b0001, 4'b1110, 4'b1000, 4'b1101, 4'b0110, 4'b0010, 4'b1011, 4'b1111, 4'b1100,
      4'b1001, 4'b0111, 4'b0011, 4'b1010, 4'b0101, 4'b0000, 4'b1111, 4'b1100, 4'b1000,
      4'b0010, 4'b0100, 4'b1001, 4'b0001, 4'b0111, 4'b0101, 4'b1011, 4'b0011, 4'b1110,
      4'b1010, 4'b0000, 4'b0110, 4'b1101, I_1);

  function automatic [3:0] MUX_v_4_64_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [3:0] input_8;
    input [3:0] input_9;
    input [3:0] input_10;
    input [3:0] input_11;
    input [3:0] input_12;
    input [3:0] input_13;
    input [3:0] input_14;
    input [3:0] input_15;
    input [3:0] input_16;
    input [3:0] input_17;
    input [3:0] input_18;
    input [3:0] input_19;
    input [3:0] input_20;
    input [3:0] input_21;
    input [3:0] input_22;
    input [3:0] input_23;
    input [3:0] input_24;
    input [3:0] input_25;
    input [3:0] input_26;
    input [3:0] input_27;
    input [3:0] input_28;
    input [3:0] input_29;
    input [3:0] input_30;
    input [3:0] input_31;
    input [3:0] input_32;
    input [3:0] input_33;
    input [3:0] input_34;
    input [3:0] input_35;
    input [3:0] input_36;
    input [3:0] input_37;
    input [3:0] input_38;
    input [3:0] input_39;
    input [3:0] input_40;
    input [3:0] input_41;
    input [3:0] input_42;
    input [3:0] input_43;
    input [3:0] input_44;
    input [3:0] input_45;
    input [3:0] input_46;
    input [3:0] input_47;
    input [3:0] input_48;
    input [3:0] input_49;
    input [3:0] input_50;
    input [3:0] input_51;
    input [3:0] input_52;
    input [3:0] input_53;
    input [3:0] input_54;
    input [3:0] input_55;
    input [3:0] input_56;
    input [3:0] input_57;
    input [3:0] input_58;
    input [3:0] input_59;
    input [3:0] input_60;
    input [3:0] input_61;
    input [3:0] input_62;
    input [3:0] input_63;
    input [5:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_4_64_2 = result;
  end
  endfunction

endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Sun Mar 21 13:06:38 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    des_check_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module des_check_core_core_fsm (
  clk, rst, fsm_output
);
  input clk;
  input rst;
  output [16:0] fsm_output;
  reg [16:0] fsm_output;


  // FSM State Type Declaration for des_check_core_core_fsm_1
  parameter
    main_C_0 = 5'd0,
    main_C_1 = 5'd1,
    main_C_2 = 5'd2,
    main_C_3 = 5'd3,
    main_C_4 = 5'd4,
    main_C_5 = 5'd5,
    main_C_6 = 5'd6,
    main_C_7 = 5'd7,
    main_C_8 = 5'd8,
    main_C_9 = 5'd9,
    main_C_10 = 5'd10,
    main_C_11 = 5'd11,
    main_C_12 = 5'd12,
    main_C_13 = 5'd13,
    main_C_14 = 5'd14,
    main_C_15 = 5'd15,
    main_C_16 = 5'd16;

  reg [4:0] state_var;
  reg [4:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : des_check_core_core_fsm_1
    case (state_var)
      main_C_1 : begin
        fsm_output = 17'b00000000000000010;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 17'b00000000000000100;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 17'b00000000000001000;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 17'b00000000000010000;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 17'b00000000000100000;
        state_var_NS = main_C_6;
      end
      main_C_6 : begin
        fsm_output = 17'b00000000001000000;
        state_var_NS = main_C_7;
      end
      main_C_7 : begin
        fsm_output = 17'b00000000010000000;
        state_var_NS = main_C_8;
      end
      main_C_8 : begin
        fsm_output = 17'b00000000100000000;
        state_var_NS = main_C_9;
      end
      main_C_9 : begin
        fsm_output = 17'b00000001000000000;
        state_var_NS = main_C_10;
      end
      main_C_10 : begin
        fsm_output = 17'b00000010000000000;
        state_var_NS = main_C_11;
      end
      main_C_11 : begin
        fsm_output = 17'b00000100000000000;
        state_var_NS = main_C_12;
      end
      main_C_12 : begin
        fsm_output = 17'b00001000000000000;
        state_var_NS = main_C_13;
      end
      main_C_13 : begin
        fsm_output = 17'b00010000000000000;
        state_var_NS = main_C_14;
      end
      main_C_14 : begin
        fsm_output = 17'b00100000000000000;
        state_var_NS = main_C_15;
      end
      main_C_15 : begin
        fsm_output = 17'b01000000000000000;
        state_var_NS = main_C_16;
      end
      main_C_16 : begin
        fsm_output = 17'b10000000000000000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 17'b00000000000000001;
        state_var_NS = main_C_1;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    des_check_core
// ------------------------------------------------------------------


module des_check_core (
  clk, rst, input_rsc_dat, input_rsc_triosy_lz, key_rsc_dat, key_rsc_triosy_lz, return_rsc_dat,
      return_rsc_triosy_lz
);
  input clk;
  input rst;
  input [63:0] input_rsc_dat;
  output input_rsc_triosy_lz;
  input [63:0] key_rsc_dat;
  output key_rsc_triosy_lz;
  output [63:0] return_rsc_dat;
  output return_rsc_triosy_lz;


  // Interconnect Declarations
  wire [63:0] input_rsci_idat;
  wire [63:0] key_rsci_idat;
  reg return_rsc_triosy_obj_ld;
  reg return_rsci_idat_63;
  reg return_rsci_idat_62;
  reg return_rsci_idat_61;
  reg return_rsci_idat_60;
  reg return_rsci_idat_59;
  reg return_rsci_idat_58;
  reg return_rsci_idat_57;
  reg return_rsci_idat_56;
  reg return_rsci_idat_55;
  reg return_rsci_idat_54;
  reg return_rsci_idat_53;
  reg return_rsci_idat_52;
  reg return_rsci_idat_51;
  reg return_rsci_idat_50;
  reg return_rsci_idat_49;
  reg return_rsci_idat_48;
  reg return_rsci_idat_47;
  reg return_rsci_idat_46;
  reg return_rsci_idat_45;
  reg return_rsci_idat_44;
  reg return_rsci_idat_43;
  reg return_rsci_idat_42;
  reg return_rsci_idat_41;
  reg return_rsci_idat_40;
  reg return_rsci_idat_39;
  reg return_rsci_idat_38;
  reg return_rsci_idat_37;
  reg return_rsci_idat_36;
  reg return_rsci_idat_35;
  reg return_rsci_idat_34;
  reg return_rsci_idat_33;
  reg return_rsci_idat_32;
  reg return_rsci_idat_31;
  reg return_rsci_idat_30;
  reg return_rsci_idat_29;
  reg return_rsci_idat_28;
  reg return_rsci_idat_27;
  reg return_rsci_idat_26;
  reg return_rsci_idat_25;
  reg return_rsci_idat_24;
  reg return_rsci_idat_23;
  reg return_rsci_idat_22;
  reg return_rsci_idat_21;
  reg return_rsci_idat_20;
  reg return_rsci_idat_19;
  reg return_rsci_idat_18;
  reg return_rsci_idat_17;
  reg return_rsci_idat_16;
  reg return_rsci_idat_15;
  reg return_rsci_idat_14;
  reg return_rsci_idat_13;
  reg return_rsci_idat_12;
  reg return_rsci_idat_11;
  reg return_rsci_idat_10;
  reg return_rsci_idat_9;
  reg return_rsci_idat_8;
  reg return_rsci_idat_7;
  reg return_rsci_idat_6;
  reg return_rsci_idat_5;
  reg return_rsci_idat_4;
  reg return_rsci_idat_3;
  reg return_rsci_idat_2;
  reg return_rsci_idat_1;
  reg return_rsci_idat_0;
  wire [16:0] fsm_output;
  reg [62:0] reg_input_ftd;
  wire R_or_1_cse;
  reg reg_key_rsc_triosy_obj_ld_cse;
  wire R_or_2_cse;
  wire R_or_8_cse;
  wire R_or_4_cse;
  wire R_or_26_cse;
  wire R_or_32_cse;
  wire R_or_38_cse;
  wire R_or_39_cse;
  wire R_or_66_cse;
  wire [3:0] O_1_out;
  wire [3:0] O_1_out_1;
  wire [3:0] O_1_out_2;
  wire [3:0] O_1_out_3;
  wire [3:0] O_1_out_4;
  wire [3:0] O_1_out_5;
  wire [3:0] O_1_out_6;
  wire [3:0] O_1_out_7;
  wire [3:0] O_1_out_8;
  reg [62:0] key_io_read_key_rsc_cse_63_1_sva;
  reg R_15_1_sva;
  reg R_11_1_sva;
  reg R_20_1_sva;
  reg R_10_1_sva;
  reg R_7_1_sva;
  reg R_3_1_sva;
  reg R_0_1_sva;
  reg [3:0] s_output_1_19_16_20_sva;
  reg [3:0] s_output_1_3_0_24_sva;
  reg [3:0] s_output_1_19_16_35_sva;
  reg [3:0] s_output_1_3_0_39_sva;
  reg [3:0] s_output_1_19_16_50_sva;
  reg [3:0] s_output_1_3_0_54_sva;
  reg [3:0] s_output_1_19_16_5_sva;
  reg [3:0] s_output_1_3_0_9_sva;
  reg R_16_3_sva;
  reg R_14_3_sva;
  reg R_18_3_sva;
  reg R_11_3_sva;
  reg R_21_3_sva;
  reg R_7_3_sva;
  reg R_24_3_sva;
  reg R_3_3_sva;
  reg R_2_3_sva;
  reg R_31_3_sva;
  reg R_15_4_sva;
  reg R_16_4_sva;
  reg R_12_4_sva;
  reg R_19_4_sva;
  reg R_11_4_sva;
  reg R_20_4_sva;
  reg R_9_4_sva;
  reg R_8_4_sva;
  reg R_23_4_sva;
  reg R_7_4_sva;
  reg R_24_4_sva;
  reg R_26_4_sva;
  reg R_4_4_sva;
  reg R_27_4_sva;
  reg R_3_4_sva;
  reg R_28_4_sva;
  reg R_29_4_sva;
  reg R_1_4_sva;
  reg R_30_4_sva;
  reg R_0_4_sva;
  reg R_31_4_sva;
  reg R_6_5_sva;
  reg R_26_5_sva;
  reg R_29_5_sva;
  reg R_25_6_sva;
  reg R_1_6_sva;
  reg R_21_7_sva;
  reg R_22_7_sva;
  reg R_1_7_sva;
  reg R_1_8_sva;
  reg R_15_9_sva;
  reg R_1_9_sva;
  reg R_0_9_sva;
  reg R_15_10_sva;
  reg R_10_10_sva;
  reg R_27_10_sva;
  reg R_0_10_sva;
  reg R_31_10_sva;
  reg R_15_11_sva;
  reg R_12_11_sva;
  reg R_19_11_sva;
  reg R_11_11_sva;
  reg R_20_11_sva;
  reg R_23_11_sva;
  reg R_7_11_sva;
  reg R_24_11_sva;
  reg R_4_11_sva;
  reg R_27_11_sva;
  reg R_3_11_sva;
  reg R_28_11_sva;
  reg R_0_11_sva;
  reg R_31_11_sva;
  reg R_1_14_sva;
  wire loop_DES_rounds_9_xor_81;
  wire loop_DES_rounds_5_xor_81;
  wire loop_DES_rounds_7_xor_81;
  wire loop_DES_rounds_8_xor_81;
  wire loop_DES_rounds_6_xor_81;
  wire loop_DES_rounds_9_xor_83;
  wire loop_DES_rounds_8_xor_83;
  wire loop_DES_rounds_10_xor_81;
  wire loop_DES_rounds_8_xor_85;
  wire loop_DES_rounds_10_xor_83;
  wire loop_DES_rounds_4_xor_81;
  wire loop_DES_rounds_7_xor_83;
  wire loop_DES_rounds_4_xor_83;
  wire loop_DES_rounds_9_xor_85;
  wire loop_DES_rounds_4_xor_85;
  wire loop_DES_rounds_8_xor_87;
  wire loop_DES_rounds_4_xor_87;
  wire loop_DES_rounds_10_xor_85;
  wire loop_DES_rounds_2_xor_81;
  wire loop_DES_rounds_10_xor_87;
  wire loop_DES_rounds_6_xor_83;
  wire loop_DES_rounds_4_xor_89;
  wire loop_DES_rounds_2_xor_83;
  wire loop_DES_rounds_2_xor_85;
  wire loop_DES_rounds_9_xor_87;
  wire loop_DES_rounds_2_xor_87;
  wire loop_DES_rounds_8_xor_89;
  wire loop_DES_rounds_5_xor_83;
  wire loop_DES_rounds_10_xor_89;
  wire loop_DES_rounds_6_xor_85;
  wire loop_DES_rounds_7_xor_85;
  wire loop_DES_rounds_9_xor_89;
  wire loop_DES_rounds_2_xor_89;
  wire loop_DES_rounds_6_xor_87;
  wire loop_DES_rounds_4_xor_91;
  wire loop_DES_rounds_7_xor_87;
  wire loop_DES_rounds_4_xor_93;
  wire loop_DES_rounds_5_xor_85;
  wire loop_DES_rounds_2_xor_91;
  wire loop_DES_rounds_5_xor_87;
  wire loop_DES_rounds_9_xor_91;
  wire loop_DES_rounds_6_xor_89;
  wire loop_DES_rounds_5_xor_89;
  wire loop_DES_rounds_14_xor_81;
  wire loop_DES_rounds_4_xor_95;
  wire loop_DES_rounds_2_xor_93;
  wire loop_DES_rounds_6_xor_91;
  wire loop_DES_rounds_4_xor_97;
  wire loop_DES_rounds_2_xor_95;
  wire loop_DES_rounds_6_xor_93;
  wire loop_DES_rounds_9_xor_93;
  wire [3:0] ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_16;
  wire [3:0] ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_17;
  wire [3:0] ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_16;
  wire [3:0] ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_16;
  wire [3:0] ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_16;
  wire [3:0] ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_16;
  wire [3:0] ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_17;
  wire [3:0] ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_17;
  wire [3:0] ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_17;
  wire [3:0] ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_17;
  wire [3:0] ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_17;
  wire [3:0] ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_17;
  wire loop_DES_rounds_16_xor_21_cse;
  wire loop_DES_rounds_16_xor_25_cse;
  wire loop_DES_rounds_16_xor_17_cse;
  wire R_or_133_cse;
  wire loop_DES_rounds_16_xor_5_cse;
  wire loop_DES_rounds_16_xor_10_cse;
  wire loop_DES_rounds_16_xor_9_cse;
  wire loop_DES_rounds_10_xor_14_cse;
  wire loop_DES_rounds_16_xor_31_cse;
  wire R_or_127_cse;
  wire R_or_120_cse;
  wire loop_DES_rounds_16_xor_4_cse;
  wire loop_DES_rounds_8_xor_4_cse;
  wire loop_DES_rounds_5_xor_1_cse;
  wire R_or_118_cse;
  wire loop_DES_rounds_16_xor_18_cse;
  wire R_or_cse;
  wire R_or_122_cse;
  wire loop_DES_rounds_16_xor_24_cse;
  wire loop_DES_rounds_16_xor_26_cse;
  wire loop_DES_rounds_16_xor_32_cse;
  wire loop_DES_rounds_16_xor_23_cse;
  wire loop_DES_rounds_11_xor_17_cse;
  wire loop_DES_rounds_5_xor_15_cse;
  wire loop_DES_rounds_3_xor_15_cse;
  wire loop_DES_rounds_6_xor_16_cse;
  wire loop_DES_rounds_4_xor_16_cse;
  wire loop_DES_rounds_11_xor_9_cse;
  wire loop_DES_rounds_11_xor_2_cse;
  wire loop_DES_rounds_5_xor_6_cse;
  wire loop_DES_rounds_11_xor_32_cse;
  wire loop_DES_rounds_16_xor_8_cse;
  wire loop_DES_rounds_5_xor_12_cse;
  wire loop_DES_rounds_11_xor_13_cse;
  wire loop_DES_rounds_13_xor_4_cse;
  wire loop_DES_rounds_3_xor_31_cse;
  wire loop_DES_rounds_10_xor_31_cse;
  wire loop_DES_rounds_4_xor_29_cse;
  wire loop_DES_rounds_15_xor_29_cse;
  wire loop_DES_rounds_11_xor_11_cse;
  wire loop_DES_rounds_10_xor_9_cse;
  wire loop_DES_rounds_16_xor_7_cse;
  wire loop_DES_rounds_9_xor_5_cse;
  wire loop_DES_rounds_5_xor_7_cse;
  wire loop_DES_rounds_10_xor_7_cse;
  wire loop_DES_rounds_11_xor_4_cse;
  wire loop_DES_rounds_3_xor_1_cse;
  wire loop_DES_rounds_10_xor_1_cse;
  wire loop_DES_rounds_16_xor_2_cse;
  wire loop_DES_rounds_10_xor_2_cse;
  wire loop_DES_rounds_10_xor_8_cse;
  wire loop_DES_rounds_16_xor_27_cse;
  wire loop_DES_rounds_10_xor_10_cse;
  wire loop_DES_rounds_16_xor_12_cse;
  wire loop_DES_rounds_11_xor_20_cse;
  wire loop_DES_rounds_5_xor_18_cse;
  wire loop_DES_rounds_10_xor_18_cse;
  wire loop_DES_rounds_16_xor_20_cse;
  wire loop_DES_rounds_6_xor_24_cse;
  wire loop_DES_rounds_10_xor_26_cse;
  wire loop_DES_rounds_16_xor_28_cse;
  wire loop_DES_rounds_5_xor_25_cse;
  wire loop_DES_rounds_10_xor_25_cse;
  wire loop_DES_rounds_16_xor_30_cse;
  wire loop_DES_rounds_6_xor_32_cse;
  wire loop_DES_rounds_5_xor_23_cse;
  wire loop_DES_rounds_10_xor_23_cse;
  wire loop_DES_rounds_6_xor_21_cse;
  wire loop_DES_rounds_10_xor_17_cse;
  wire loop_DES_rounds_16_xor_15_cse;
  wire loop_DES_rounds_10_xor_15_cse;
  wire loop_DES_rounds_5_xor_11_cse;
  wire loop_DES_rounds_5_xor_29_cse;
  wire loop_DES_rounds_6_xor_6_cse;
  wire loop_DES_rounds_4_xor_3_cse;
  wire loop_DES_rounds_5_xor_27_cse;
  wire loop_DES_rounds_16_xor_14_cse;
  wire loop_DES_rounds_11_xor_12_cse;
  wire loop_DES_rounds_10_xor_20_cse;
  wire loop_DES_rounds_16_xor_22_cse;
  wire loop_DES_rounds_5_xor_30_cse;
  wire R_or_105_cse;
  wire loop_DES_rounds_13_xor_13_cse;
  wire loop_DES_rounds_13_xor_19_cse;
  wire loop_DES_rounds_11_xor_19_cse;
  wire loop_DES_rounds_10_xor_30_cse;
  wire loop_DES_rounds_6_xor_19_cse;
  wire loop_DES_rounds_16_xor_19_cse;
  wire loop_DES_rounds_10_xor_28_cse;
  wire loop_DES_rounds_5_xor_21_cse;
  wire loop_DES_rounds_15_xor_21_cse;
  wire loop_DES_rounds_10_xor_22_cse;
  wire loop_DES_rounds_7_xor_28_cse;
  wire loop_DES_rounds_15_xor_28_cse;
  wire loop_DES_rounds_13_xor_30_cse;
  wire loop_DES_rounds_12_xor_13_cse;
  wire loop_DES_rounds_10_xor_13_cse;
  wire loop_DES_rounds_11_xor_14_cse;
  wire loop_DES_rounds_7_xor_22_cse;

  wire[0:0] loop_DES_rounds_1_xor_31_nl;
  wire[0:0] loop_DES_rounds_2_xor_31_nl;
  wire[0:0] loop_DES_rounds_15_xor_3_nl;
  wire[0:0] loop_DES_rounds_1_xor_25_nl;
  wire[0:0] loop_DES_rounds_2_xor_25_nl;
  wire[0:0] loop_DES_rounds_8_xor_5_nl;
  wire[0:0] loop_DES_rounds_1_xor_17_nl;
  wire[0:0] loop_DES_rounds_2_xor_17_nl;
  wire[0:0] loop_DES_rounds_5_xor_3_nl;
  wire[0:0] loop_DES_rounds_7_xor_6_nl;
  wire[0:0] loop_DES_rounds_1_xor_11_nl;
  wire[0:0] loop_DES_rounds_2_xor_19_nl;
  wire[0:0] loop_DES_rounds_8_xor_11_nl;
  wire[0:0] loop_DES_rounds_12_xor_6_nl;
  wire[0:0] loop_DES_rounds_14_xor_3_nl;
  wire[0:0] loop_DES_rounds_1_xor_10_nl;
  wire[0:0] loop_DES_rounds_2_xor_10_nl;
  wire[0:0] loop_DES_rounds_6_xor_27_nl;
  wire[0:0] loop_DES_rounds_1_xor_9_nl;
  wire[0:0] loop_DES_rounds_2_xor_9_nl;
  wire[0:0] loop_DES_rounds_4_xor_14_nl;
  wire[0:0] loop_DES_rounds_7_xor_27_nl;
  wire[0:0] loop_DES_rounds_1_xor_1_nl;
  wire[0:0] loop_DES_rounds_2_xor_1_nl;
  wire[0:0] loop_DES_rounds_6_xor_14_nl;
  wire[0:0] loop_DES_rounds_13_xor_20_nl;
  wire[0:0] loop_DES_rounds_1_xor_29_nl;
  wire[0:0] loop_DES_rounds_1_xor_5_nl;
  wire[0:0] loop_DES_rounds_3_xor_7_nl;
  wire[0:0] loop_DES_rounds_13_xor_9_nl;
  wire[0:0] loop_DES_rounds_1_xor_2_nl;
  wire[0:0] loop_DES_rounds_1_xor_16_nl;
  wire[0:0] loop_DES_rounds_13_xor_2_nl;
  wire[0:0] loop_DES_rounds_1_xor_27_nl;
  wire[0:0] loop_DES_rounds_3_xor_8_nl;
  wire[0:0] loop_DES_rounds_5_xor_8_nl;
  wire[0:0] loop_DES_rounds_1_xor_12_nl;
  wire[0:0] loop_DES_rounds_5_xor_10_nl;
  wire[0:0] loop_DES_rounds_1_xor_18_nl;
  wire[0:0] loop_DES_rounds_3_xor_16_nl;
  wire[0:0] loop_DES_rounds_5_xor_16_nl;
  wire[0:0] loop_DES_rounds_1_xor_4_nl;
  wire[0:0] loop_DES_rounds_2_xor_18_nl;
  wire[0:0] loop_DES_rounds_1_xor_20_nl;
  wire[0:0] loop_DES_rounds_3_xor_18_nl;
  wire[0:0] loop_DES_rounds_11_xor_5_nl;
  wire[0:0] loop_DES_rounds_13_xor_6_nl;
  wire[0:0] loop_DES_rounds_1_xor_26_nl;
  wire[0:0] loop_DES_rounds_3_xor_24_nl;
  wire[0:0] loop_DES_rounds_5_xor_24_nl;
  wire[0:0] loop_DES_rounds_1_xor_6_nl;
  wire[0:0] loop_DES_rounds_2_xor_26_nl;
  wire[0:0] loop_DES_rounds_1_xor_28_nl;
  wire[0:0] loop_DES_rounds_3_xor_26_nl;
  wire[0:0] loop_DES_rounds_5_xor_26_nl;
  wire[0:0] loop_DES_rounds_1_xor_21_nl;
  wire[0:0] loop_DES_rounds_3_xor_23_nl;
  wire[0:0] loop_DES_rounds_13_xor_32_nl;
  wire[0:0] loop_DES_rounds_1_xor_24_nl;
  wire[0:0] loop_DES_rounds_2_xor_23_nl;
  wire[0:0] loop_DES_rounds_1_xor_13_nl;
  wire[0:0] loop_DES_rounds_13_xor_17_nl;
  wire[0:0] loop_DES_rounds_1_xor_15_nl;
  wire[0:0] loop_DES_rounds_1_xor_22_nl;
  wire[0:0] loop_DES_rounds_2_xor_16_nl;
  wire[0:0] loop_DES_rounds_8_xor_29_nl;
  wire[0:0] loop_DES_rounds_1_xor_3_nl;
  wire[0:0] loop_DES_rounds_3_xor_29_nl;
  wire[0:0] loop_DES_rounds_7_xor_11_nl;
  wire[0:0] loop_DES_rounds_11_xor_31_nl;
  wire[0:0] loop_DES_rounds_13_xor_31_nl;
  wire[0:0] loop_DES_rounds_1_xor_7_nl;
  wire[0:0] loop_DES_rounds_15_xor_5_nl;
  wire[0:0] loop_DES_rounds_1_xor_8_nl;
  wire[0:0] loop_DES_rounds_3_xor_2_nl;
  wire[0:0] loop_DES_rounds_1_xor_30_nl;
  wire[0:0] loop_DES_rounds_13_xor_5_nl;
  wire[0:0] loop_DES_rounds_1_xor_23_nl;
  wire[0:0] loop_DES_rounds_3_xor_32_nl;
  wire[0:0] loop_DES_rounds_11_xor_3_nl;
  wire[0:0] loop_DES_rounds_14_xor_6_nl;
  wire[0:0] loop_DES_rounds_1_xor_19_nl;
  wire[0:0] loop_DES_rounds_2_xor_6_nl;
  wire[0:0] loop_DES_rounds_6_xor_3_nl;
  wire[0:0] loop_DES_rounds_9_xor_11_nl;
  wire[0:0] loop_DES_rounds_15_xor_6_nl;
  wire[0:0] R_or_125_nl;
  wire[0:0] loop_DES_rounds_1_xor_14_nl;
  wire[0:0] loop_DES_rounds_2_xor_8_nl;
  wire[0:0] loop_DES_rounds_4_xor_11_nl;
  wire[0:0] loop_DES_rounds_6_xor_29_nl;
  wire[0:0] loop_DES_rounds_8_xor_3_nl;
  wire[0:0] loop_DES_rounds_1_xor_32_nl;
  wire[0:0] loop_DES_rounds_3_xor_11_nl;
  wire[0:0] loop_DES_rounds_7_xor_3_nl;
  wire[0:0] loop_DES_rounds_13_xor_27_nl;
  wire[0:0] R_or_102_nl;
  wire[0:0] loop_DES_rounds_3_xor_27_nl;
  wire[0:0] loop_DES_rounds_9_xor_27_nl;
  wire[0:0] loop_DES_rounds_13_xor_12_nl;
  wire[0:0] loop_DES_rounds_3_xor_12_nl;
  wire[0:0] loop_DES_rounds_6_xor_12_nl;
  wire[0:0] loop_DES_rounds_13_xor_14_nl;
  wire[0:0] loop_DES_rounds_3_xor_6_nl;
  wire[0:0] loop_DES_rounds_9_xor_6_nl;
  wire[0:0] loop_DES_rounds_15_xor_27_nl;
  wire[0:0] loop_DES_rounds_3_xor_3_nl;
  wire[0:0] loop_DES_rounds_5_xor_13_nl;
  wire[0:0] loop_DES_rounds_2_xor_29_nl;
  wire[0:0] loop_DES_rounds_10_xor_29_nl;
  wire[0:0] loop_DES_rounds_2_xor_11_nl;
  wire[0:0] loop_DES_rounds_11_xor_29_nl;
  wire[0:0] loop_DES_rounds_2_xor_7_nl;
  wire[0:0] loop_DES_rounds_3_xor_5_nl;
  wire[0:0] loop_DES_rounds_9_xor_3_nl;
  wire[0:0] loop_DES_rounds_13_xor_7_nl;
  wire[0:0] R_or_99_nl;
  wire[0:0] loop_DES_rounds_2_xor_5_nl;
  wire[0:0] loop_DES_rounds_10_xor_5_nl;
  wire[0:0] loop_DES_rounds_3_xor_4_nl;
  wire[0:0] loop_DES_rounds_11_xor_1_nl;
  wire[0:0] loop_DES_rounds_13_xor_1_nl;
  wire[0:0] loop_DES_rounds_2_xor_2_nl;
  wire[0:0] loop_DES_rounds_2_xor_4_nl;
  wire[0:0] loop_DES_rounds_10_xor_4_nl;
  wire[0:0] loop_DES_rounds_2_xor_27_nl;
  wire[0:0] loop_DES_rounds_10_xor_27_nl;
  wire[0:0] loop_DES_rounds_2_xor_12_nl;
  wire[0:0] loop_DES_rounds_3_xor_20_nl;
  wire[0:0] loop_DES_rounds_13_xor_18_nl;
  wire[0:0] loop_DES_rounds_2_xor_20_nl;
  wire[0:0] loop_DES_rounds_2_xor_24_nl;
  wire[0:0] loop_DES_rounds_4_xor_6_nl;
  wire[0:0] loop_DES_rounds_6_xor_5_nl;
  wire[0:0] loop_DES_rounds_8_xor_6_nl;
  wire[0:0] loop_DES_rounds_2_xor_28_nl;
  wire[0:0] loop_DES_rounds_3_xor_30_nl;
  wire[0:0] loop_DES_rounds_13_xor_25_nl;
  wire[0:0] loop_DES_rounds_2_xor_30_nl;
  wire[0:0] loop_DES_rounds_2_xor_32_nl;
  wire[0:0] loop_DES_rounds_8_xor_27_nl;
  wire[0:0] loop_DES_rounds_3_xor_21_nl;
  wire[0:0] loop_DES_rounds_13_xor_23_nl;
  wire[0:0] loop_DES_rounds_2_xor_21_nl;
  wire[0:0] loop_DES_rounds_2_xor_15_nl;
  wire[0:0] loop_DES_rounds_2_xor_13_nl;
  wire[0:0] loop_DES_rounds_2_xor_3_nl;
  wire[0:0] loop_DES_rounds_4_xor_19_nl;
  wire[0:0] loop_DES_rounds_10_xor_3_nl;
  wire[0:0] loop_DES_rounds_2_xor_14_nl;
  wire[0:0] loop_DES_rounds_14_xor_11_nl;
  wire[0:0] loop_DES_rounds_2_xor_22_nl;
  wire[0:0] loop_DES_rounds_6_xor_11_nl;
  wire[0:0] loop_DES_rounds_9_xor_29_nl;
  wire[0:0] loop_DES_rounds_13_xor_3_nl;
  wire[0:0] loop_DES_rounds_3_xor_14_nl;
  wire[0:0] loop_DES_rounds_7_xor_12_nl;
  wire[0:0] loop_DES_rounds_12_xor_14_nl;
  wire[0:0] R_or_152_nl;
  wire[0:0] loop_DES_rounds_3_xor_22_nl;
  wire[0:0] loop_DES_rounds_6_xor_20_nl;
  wire[0:0] loop_DES_rounds_3_xor_28_nl;
  wire[0:0] loop_DES_rounds_3_xor_19_nl;
  wire[0:0] loop_DES_rounds_5_xor_28_nl;
  wire[0:0] loop_DES_rounds_3_xor_13_nl;
  wire[0:0] loop_DES_rounds_4_xor_22_nl;
  wire[0:0] loop_DES_rounds_13_xor_22_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [63:0] nl_return_rsci_idat;
  assign nl_return_rsci_idat = {return_rsci_idat_63 , return_rsci_idat_62 , return_rsci_idat_61
      , return_rsci_idat_60 , return_rsci_idat_59 , return_rsci_idat_58 , return_rsci_idat_57
      , return_rsci_idat_56 , return_rsci_idat_55 , return_rsci_idat_54 , return_rsci_idat_53
      , return_rsci_idat_52 , return_rsci_idat_51 , return_rsci_idat_50 , return_rsci_idat_49
      , return_rsci_idat_48 , return_rsci_idat_47 , return_rsci_idat_46 , return_rsci_idat_45
      , return_rsci_idat_44 , return_rsci_idat_43 , return_rsci_idat_42 , return_rsci_idat_41
      , return_rsci_idat_40 , return_rsci_idat_39 , return_rsci_idat_38 , return_rsci_idat_37
      , return_rsci_idat_36 , return_rsci_idat_35 , return_rsci_idat_34 , return_rsci_idat_33
      , return_rsci_idat_32 , return_rsci_idat_31 , return_rsci_idat_30 , return_rsci_idat_29
      , return_rsci_idat_28 , return_rsci_idat_27 , return_rsci_idat_26 , return_rsci_idat_25
      , return_rsci_idat_24 , return_rsci_idat_23 , return_rsci_idat_22 , return_rsci_idat_21
      , return_rsci_idat_20 , return_rsci_idat_19 , return_rsci_idat_18 , return_rsci_idat_17
      , return_rsci_idat_16 , return_rsci_idat_15 , return_rsci_idat_14 , return_rsci_idat_13
      , return_rsci_idat_12 , return_rsci_idat_11 , return_rsci_idat_10 , return_rsci_idat_9
      , return_rsci_idat_8 , return_rsci_idat_7 , return_rsci_idat_6 , return_rsci_idat_5
      , return_rsci_idat_4 , return_rsci_idat_3 , return_rsci_idat_2 , return_rsci_idat_1
      , return_rsci_idat_0};
  wire[0:0] loop_DES_rounds_xor_nl;
  wire[0:0] loop_DES_rounds_xor_1_nl;
  wire[0:0] loop_DES_rounds_xor_2_nl;
  wire[0:0] loop_DES_rounds_xor_3_nl;
  wire[0:0] loop_DES_rounds_xor_4_nl;
  wire[0:0] loop_DES_rounds_xor_5_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_1_rg_I_1;
  assign loop_DES_rounds_xor_nl = (input_rsci_idat[30]) ^ (ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_17[3])
      ^ (key_rsci_idat[39]);
  assign loop_DES_rounds_xor_1_nl = (input_rsci_idat[4]) ^ (O_1_out_3[3]) ^ (key_rsci_idat[30]);
  assign loop_DES_rounds_xor_2_nl = (input_rsci_idat[38]) ^ (ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_17[3])
      ^ (key_rsci_idat[15]);
  assign loop_DES_rounds_xor_3_nl = (input_rsci_idat[46]) ^ (ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_17[0])
      ^ (key_rsci_idat[5]);
  assign loop_DES_rounds_xor_4_nl = (input_rsci_idat[54]) ^ (ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_17[0])
      ^ (key_rsci_idat[63]);
  assign loop_DES_rounds_xor_5_nl = (input_rsci_idat[62]) ^ (ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_17[3])
      ^ (key_rsci_idat[53]);
  assign nl_U_ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_1_rg_I_1 = {loop_DES_rounds_xor_nl
      , loop_DES_rounds_xor_1_nl , loop_DES_rounds_xor_2_nl , loop_DES_rounds_xor_3_nl
      , loop_DES_rounds_xor_4_nl , loop_DES_rounds_xor_5_nl};
  wire[0:0] loop_DES_rounds_2_xor_50_nl;
  wire[0:0] loop_DES_rounds_2_xor_55_nl;
  wire[0:0] loop_DES_rounds_xor_8_nl;
  wire[0:0] loop_DES_rounds_2_xor_52_nl;
  wire[0:0] loop_DES_rounds_2_xor_54_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_1_rg_I_1;
  assign loop_DES_rounds_2_xor_50_nl = R_20_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_2_xor_55_nl = R_15_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign loop_DES_rounds_xor_8_nl = (reg_input_ftd[35]) ^ (ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_17[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_2_xor_52_nl = R_27_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_2_xor_54_nl = R_15_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign nl_U_ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_1_rg_I_1 = {loop_DES_rounds_2_xor_50_nl
      , loop_DES_rounds_2_xor_55_nl , loop_DES_rounds_xor_8_nl , loop_DES_rounds_2_xor_52_nl
      , loop_DES_rounds_2_xor_81 , loop_DES_rounds_2_xor_54_nl};
  wire[0:0] loop_DES_rounds_2_xor_68_nl;
  wire[0:0] loop_DES_rounds_2_xor_73_nl;
  wire[0:0] loop_DES_rounds_2_xor_69_nl;
  wire[0:0] loop_DES_rounds_xor_9_nl;
  wire[0:0] loop_DES_rounds_2_xor_71_nl;
  wire[0:0] loop_DES_rounds_xor_10_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_1_rg_I_1;
  assign loop_DES_rounds_2_xor_68_nl = R_7_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_2_xor_73_nl = R_3_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_2_xor_69_nl = R_7_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_xor_9_nl = (reg_input_ftd[7]) ^ (s_output_1_19_16_20_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_2_xor_71_nl = R_31_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_xor_10_nl = (reg_input_ftd[23]) ^ (ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_17[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign nl_U_ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_1_rg_I_1 = {loop_DES_rounds_2_xor_68_nl
      , loop_DES_rounds_2_xor_73_nl , loop_DES_rounds_2_xor_69_nl , loop_DES_rounds_xor_9_nl
      , loop_DES_rounds_2_xor_71_nl , loop_DES_rounds_xor_10_nl};
  wire[0:0] loop_DES_rounds_2_xor_61_nl;
  wire[0:0] loop_DES_rounds_2_xor_57_nl;
  wire[0:0] loop_DES_rounds_xor_14_nl;
  wire[0:0] loop_DES_rounds_2_xor_59_nl;
  wire[0:0] loop_DES_rounds_xor_15_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_1_rg_I_1;
  assign loop_DES_rounds_2_xor_61_nl = R_11_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_2_xor_57_nl = R_15_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_xor_14_nl = (reg_input_ftd[9]) ^ (ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_17[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_2_xor_59_nl = R_11_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_xor_15_nl = (reg_input_ftd[25]) ^ (s_output_1_19_16_20_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign nl_U_ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_1_rg_I_1 = {loop_DES_rounds_2_xor_87
      , loop_DES_rounds_2_xor_61_nl , loop_DES_rounds_2_xor_57_nl , loop_DES_rounds_xor_14_nl
      , loop_DES_rounds_2_xor_59_nl , loop_DES_rounds_xor_15_nl};
  wire[0:0] loop_DES_rounds_xor_11_nl;
  wire[0:0] loop_DES_rounds_2_xor_45_nl;
  wire[0:0] loop_DES_rounds_xor_12_nl;
  wire[0:0] loop_DES_rounds_2_xor_47_nl;
  wire[0:0] loop_DES_rounds_2_xor_48_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_1_rg_I_1;
  assign loop_DES_rounds_xor_11_nl = (reg_input_ftd[35]) ^ (ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_17[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_2_xor_45_nl = R_15_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_xor_12_nl = (reg_input_ftd[11]) ^ (s_output_1_19_16_20_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_2_xor_47_nl = R_20_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_2_xor_48_nl = R_20_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign nl_U_ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_1_rg_I_1 = {loop_DES_rounds_2_xor_83
      , loop_DES_rounds_xor_11_nl , loop_DES_rounds_2_xor_45_nl , loop_DES_rounds_xor_12_nl
      , loop_DES_rounds_2_xor_47_nl , loop_DES_rounds_2_xor_48_nl};
  wire[0:0] loop_DES_rounds_xor_6_nl;
  wire[0:0] loop_DES_rounds_xor_7_nl;
  wire[0:0] loop_DES_rounds_2_xor_76_nl;
  wire[0:0] loop_DES_rounds_2_xor_77_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_1_rg_I_1;
  assign loop_DES_rounds_xor_6_nl = (reg_input_ftd[23]) ^ (ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_17[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_xor_7_nl = (reg_input_ftd[5]) ^ (s_output_1_19_16_20_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_2_xor_76_nl = R_19_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_2_xor_77_nl = R_0_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign nl_U_ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_1_rg_I_1 = {loop_DES_rounds_xor_6_nl
      , loop_DES_rounds_xor_7_nl , loop_DES_rounds_2_xor_91 , loop_DES_rounds_2_xor_76_nl
      , loop_DES_rounds_2_xor_77_nl , loop_DES_rounds_2_xor_93};
  wire[0:0] loop_DES_rounds_1_xor_74_nl;
  wire[0:0] loop_DES_rounds_1_xor_79_nl;
  wire[0:0] loop_DES_rounds_1_xor_75_nl;
  wire[0:0] loop_DES_rounds_1_xor_76_nl;
  wire[0:0] loop_DES_rounds_1_xor_77_nl;
  wire[0:0] loop_DES_rounds_1_xor_78_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_rg_I_1;
  assign loop_DES_rounds_1_xor_74_nl = (input_rsci_idat[25]) ^ (key_rsci_idat[19]);
  assign loop_DES_rounds_1_xor_79_nl = (input_rsci_idat[7]) ^ (key_rsci_idat[33]);
  assign loop_DES_rounds_1_xor_75_nl = (input_rsci_idat[33]) ^ (key_rsci_idat[50]);
  assign loop_DES_rounds_1_xor_76_nl = (input_rsci_idat[41]) ^ (key_rsci_idat[51]);
  assign loop_DES_rounds_1_xor_77_nl = (input_rsci_idat[49]) ^ (key_rsci_idat[2]);
  assign loop_DES_rounds_1_xor_78_nl = (input_rsci_idat[57]) ^ (key_rsci_idat[9]);
  assign nl_U_ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_rg_I_1 = {loop_DES_rounds_1_xor_74_nl
      , loop_DES_rounds_1_xor_79_nl , loop_DES_rounds_1_xor_75_nl , loop_DES_rounds_1_xor_76_nl
      , loop_DES_rounds_1_xor_77_nl , loop_DES_rounds_1_xor_78_nl};
  wire[0:0] loop_DES_rounds_1_xor_68_nl;
  wire[0:0] loop_DES_rounds_1_xor_73_nl;
  wire[0:0] loop_DES_rounds_1_xor_69_nl;
  wire[0:0] loop_DES_rounds_1_xor_70_nl;
  wire[0:0] loop_DES_rounds_1_xor_71_nl;
  wire[0:0] loop_DES_rounds_1_xor_72_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_rg_I_1;
  assign loop_DES_rounds_1_xor_68_nl = (input_rsci_idat[59]) ^ (key_rsci_idat[3]);
  assign loop_DES_rounds_1_xor_73_nl = (input_rsci_idat[33]) ^ (key_rsci_idat[44]);
  assign loop_DES_rounds_1_xor_69_nl = (input_rsci_idat[1]) ^ (key_rsci_idat[43]);
  assign loop_DES_rounds_1_xor_70_nl = (input_rsci_idat[9]) ^ (key_rsci_idat[26]);
  assign loop_DES_rounds_1_xor_71_nl = (input_rsci_idat[17]) ^ (key_rsci_idat[1]);
  assign loop_DES_rounds_1_xor_72_nl = (input_rsci_idat[25]) ^ (key_rsci_idat[49]);
  assign nl_U_ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_rg_I_1 = {loop_DES_rounds_1_xor_68_nl
      , loop_DES_rounds_1_xor_73_nl , loop_DES_rounds_1_xor_69_nl , loop_DES_rounds_1_xor_70_nl
      , loop_DES_rounds_1_xor_71_nl , loop_DES_rounds_1_xor_72_nl};
  wire[0:0] loop_DES_rounds_1_xor_44_nl;
  wire[0:0] loop_DES_rounds_1_xor_49_nl;
  wire[0:0] loop_DES_rounds_1_xor_45_nl;
  wire[0:0] loop_DES_rounds_1_xor_46_nl;
  wire[0:0] loop_DES_rounds_1_xor_47_nl;
  wire[0:0] loop_DES_rounds_1_xor_48_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_rg_I_1;
  assign loop_DES_rounds_1_xor_44_nl = (input_rsci_idat[63]) ^ (key_rsci_idat[61]);
  assign loop_DES_rounds_1_xor_49_nl = (input_rsci_idat[37]) ^ (key_rsci_idat[6]);
  assign loop_DES_rounds_1_xor_45_nl = (input_rsci_idat[5]) ^ (key_rsci_idat[29]);
  assign loop_DES_rounds_1_xor_46_nl = (input_rsci_idat[13]) ^ (key_rsci_idat[38]);
  assign loop_DES_rounds_1_xor_47_nl = (input_rsci_idat[21]) ^ (key_rsci_idat[39]);
  assign loop_DES_rounds_1_xor_48_nl = (input_rsci_idat[29]) ^ (key_rsci_idat[20]);
  assign nl_U_ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_rg_I_1 = {loop_DES_rounds_1_xor_44_nl
      , loop_DES_rounds_1_xor_49_nl , loop_DES_rounds_1_xor_45_nl , loop_DES_rounds_1_xor_46_nl
      , loop_DES_rounds_1_xor_47_nl , loop_DES_rounds_1_xor_48_nl};
  wire[0:0] loop_DES_rounds_1_xor_62_nl;
  wire[0:0] loop_DES_rounds_1_xor_67_nl;
  wire[0:0] loop_DES_rounds_1_xor_63_nl;
  wire[0:0] loop_DES_rounds_1_xor_64_nl;
  wire[0:0] loop_DES_rounds_1_xor_65_nl;
  wire[0:0] loop_DES_rounds_1_xor_66_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_rg_I_1;
  assign loop_DES_rounds_1_xor_62_nl = (input_rsci_idat[27]) ^ (key_rsci_idat[17]);
  assign loop_DES_rounds_1_xor_67_nl = (input_rsci_idat[1]) ^ (key_rsci_idat[35]);
  assign loop_DES_rounds_1_xor_63_nl = (input_rsci_idat[35]) ^ (key_rsci_idat[34]);
  assign loop_DES_rounds_1_xor_64_nl = (input_rsci_idat[43]) ^ (key_rsci_idat[59]);
  assign loop_DES_rounds_1_xor_65_nl = (input_rsci_idat[51]) ^ (key_rsci_idat[11]);
  assign loop_DES_rounds_1_xor_66_nl = (input_rsci_idat[59]) ^ (key_rsci_idat[41]);
  assign nl_U_ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_rg_I_1 = {loop_DES_rounds_1_xor_62_nl
      , loop_DES_rounds_1_xor_67_nl , loop_DES_rounds_1_xor_63_nl , loop_DES_rounds_1_xor_64_nl
      , loop_DES_rounds_1_xor_65_nl , loop_DES_rounds_1_xor_66_nl};
  wire[0:0] loop_DES_rounds_1_xor_56_nl;
  wire[0:0] loop_DES_rounds_1_xor_61_nl;
  wire[0:0] loop_DES_rounds_1_xor_57_nl;
  wire[0:0] loop_DES_rounds_1_xor_58_nl;
  wire[0:0] loop_DES_rounds_1_xor_59_nl;
  wire[0:0] loop_DES_rounds_1_xor_60_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_rg_I_1;
  assign loop_DES_rounds_1_xor_56_nl = (input_rsci_idat[61]) ^ (key_rsci_idat[42]);
  assign loop_DES_rounds_1_xor_61_nl = (input_rsci_idat[35]) ^ (key_rsci_idat[60]);
  assign loop_DES_rounds_1_xor_57_nl = (input_rsci_idat[3]) ^ (key_rsci_idat[36]);
  assign loop_DES_rounds_1_xor_58_nl = (input_rsci_idat[11]) ^ (key_rsci_idat[25]);
  assign loop_DES_rounds_1_xor_59_nl = (input_rsci_idat[19]) ^ (key_rsci_idat[10]);
  assign loop_DES_rounds_1_xor_60_nl = (input_rsci_idat[27]) ^ (key_rsci_idat[27]);
  assign nl_U_ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_rg_I_1 = {loop_DES_rounds_1_xor_56_nl
      , loop_DES_rounds_1_xor_61_nl , loop_DES_rounds_1_xor_57_nl , loop_DES_rounds_1_xor_58_nl
      , loop_DES_rounds_1_xor_59_nl , loop_DES_rounds_1_xor_60_nl};
  wire[0:0] loop_DES_rounds_1_xor_38_nl;
  wire[0:0] loop_DES_rounds_1_xor_43_nl;
  wire[0:0] loop_DES_rounds_1_xor_39_nl;
  wire[0:0] loop_DES_rounds_1_xor_40_nl;
  wire[0:0] loop_DES_rounds_1_xor_41_nl;
  wire[0:0] loop_DES_rounds_1_xor_42_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_rg_I_1;
  assign loop_DES_rounds_1_xor_38_nl = (reg_input_ftd[30]) ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign loop_DES_rounds_1_xor_43_nl = (reg_input_ftd[4]) ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign loop_DES_rounds_1_xor_39_nl = (reg_input_ftd[38]) ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_1_xor_40_nl = (reg_input_ftd[46]) ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_1_xor_41_nl = (reg_input_ftd[54]) ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_1_xor_42_nl = (reg_input_ftd[62]) ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign nl_U_ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_rg_I_1 = {loop_DES_rounds_1_xor_38_nl
      , loop_DES_rounds_1_xor_43_nl , loop_DES_rounds_1_xor_39_nl , loop_DES_rounds_1_xor_40_nl
      , loop_DES_rounds_1_xor_41_nl , loop_DES_rounds_1_xor_42_nl};
  wire[0:0] operator_8_false_1_mux1h_nl;
  wire[0:0] loop_DES_rounds_xor_48_nl;
  wire[0:0] loop_DES_rounds_4_xor_38_nl;
  wire[0:0] loop_DES_rounds_5_xor_38_nl;
  wire[0:0] loop_DES_rounds_6_xor_38_nl;
  wire[0:0] loop_DES_rounds_8_xor_38_nl;
  wire[0:0] loop_DES_rounds_9_xor_38_nl;
  wire[0:0] loop_DES_rounds_10_xor_38_nl;
  wire[0:0] loop_DES_rounds_11_xor_38_nl;
  wire[0:0] loop_DES_rounds_12_xor_38_nl;
  wire[0:0] loop_DES_rounds_13_xor_38_nl;
  wire[0:0] loop_DES_rounds_14_xor_38_nl;
  wire[0:0] loop_DES_rounds_15_xor_38_nl;
  wire[0:0] loop_DES_rounds_16_xor_38_nl;
  wire[0:0] operator_8_false_1_mux1h_8_nl;
  wire[0:0] loop_DES_rounds_xor_49_nl;
  wire[0:0] loop_DES_rounds_6_xor_43_nl;
  wire[0:0] loop_DES_rounds_8_xor_43_nl;
  wire[0:0] loop_DES_rounds_9_xor_43_nl;
  wire[0:0] loop_DES_rounds_10_xor_43_nl;
  wire[0:0] loop_DES_rounds_11_xor_43_nl;
  wire[0:0] loop_DES_rounds_12_xor_43_nl;
  wire[0:0] loop_DES_rounds_13_xor_43_nl;
  wire[0:0] loop_DES_rounds_14_xor_43_nl;
  wire[0:0] loop_DES_rounds_15_xor_43_nl;
  wire[0:0] loop_DES_rounds_16_xor_43_nl;
  wire[0:0] operator_8_false_1_mux1h_9_nl;
  wire[0:0] loop_DES_rounds_xor_50_nl;
  wire[0:0] loop_DES_rounds_4_xor_39_nl;
  wire[0:0] loop_DES_rounds_5_xor_39_nl;
  wire[0:0] loop_DES_rounds_6_xor_39_nl;
  wire[0:0] loop_DES_rounds_7_xor_39_nl;
  wire[0:0] loop_DES_rounds_8_xor_39_nl;
  wire[0:0] loop_DES_rounds_9_xor_39_nl;
  wire[0:0] loop_DES_rounds_10_xor_39_nl;
  wire[0:0] loop_DES_rounds_11_xor_39_nl;
  wire[0:0] loop_DES_rounds_12_xor_39_nl;
  wire[0:0] loop_DES_rounds_13_xor_39_nl;
  wire[0:0] loop_DES_rounds_14_xor_39_nl;
  wire[0:0] loop_DES_rounds_15_xor_39_nl;
  wire[0:0] loop_DES_rounds_16_xor_39_nl;
  wire[0:0] operator_8_false_1_mux1h_10_nl;
  wire[0:0] loop_DES_rounds_xor_51_nl;
  wire[0:0] loop_DES_rounds_5_xor_40_nl;
  wire[0:0] loop_DES_rounds_6_xor_40_nl;
  wire[0:0] loop_DES_rounds_7_xor_40_nl;
  wire[0:0] loop_DES_rounds_8_xor_40_nl;
  wire[0:0] loop_DES_rounds_9_xor_40_nl;
  wire[0:0] loop_DES_rounds_11_xor_40_nl;
  wire[0:0] loop_DES_rounds_12_xor_40_nl;
  wire[0:0] loop_DES_rounds_13_xor_40_nl;
  wire[0:0] loop_DES_rounds_14_xor_40_nl;
  wire[0:0] loop_DES_rounds_15_xor_40_nl;
  wire[0:0] loop_DES_rounds_16_xor_40_nl;
  wire[0:0] operator_8_false_1_mux1h_11_nl;
  wire[0:0] loop_DES_rounds_xor_52_nl;
  wire[0:0] loop_DES_rounds_4_xor_41_nl;
  wire[0:0] loop_DES_rounds_5_xor_41_nl;
  wire[0:0] loop_DES_rounds_7_xor_41_nl;
  wire[0:0] loop_DES_rounds_11_xor_41_nl;
  wire[0:0] loop_DES_rounds_14_xor_41_nl;
  wire[0:0] loop_DES_rounds_16_xor_41_nl;
  wire[0:0] operator_8_false_1_mux1h_12_nl;
  wire[0:0] loop_DES_rounds_xor_53_nl;
  wire[0:0] loop_DES_rounds_4_xor_42_nl;
  wire[0:0] loop_DES_rounds_6_xor_42_nl;
  wire[0:0] loop_DES_rounds_8_xor_42_nl;
  wire[0:0] loop_DES_rounds_9_xor_42_nl;
  wire[0:0] loop_DES_rounds_10_xor_42_nl;
  wire[0:0] loop_DES_rounds_11_xor_42_nl;
  wire[0:0] loop_DES_rounds_12_xor_42_nl;
  wire[0:0] loop_DES_rounds_13_xor_42_nl;
  wire[0:0] loop_DES_rounds_14_xor_42_nl;
  wire[0:0] loop_DES_rounds_15_xor_42_nl;
  wire[0:0] loop_DES_rounds_16_xor_42_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_10_rg_I_1;
  assign loop_DES_rounds_xor_48_nl = (key_io_read_key_rsc_cse_63_1_sva[54]) ^ (reg_input_ftd[30])
      ^ (s_output_1_3_0_39_sva[3]);
  assign loop_DES_rounds_4_xor_38_nl = R_28_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_5_xor_38_nl = R_28_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign loop_DES_rounds_6_xor_38_nl = R_28_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign loop_DES_rounds_8_xor_38_nl = R_28_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign loop_DES_rounds_9_xor_38_nl = R_28_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_10_xor_38_nl = R_28_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign loop_DES_rounds_11_xor_38_nl = R_27_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_12_xor_38_nl = R_28_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_13_xor_38_nl = R_27_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_14_xor_38_nl = R_28_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign loop_DES_rounds_15_xor_38_nl = R_27_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign loop_DES_rounds_16_xor_38_nl = R_28_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign operator_8_false_1_mux1h_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_48_nl,
      loop_DES_rounds_4_xor_38_nl, loop_DES_rounds_5_xor_38_nl, loop_DES_rounds_6_xor_38_nl,
      loop_DES_rounds_7_xor_85, loop_DES_rounds_8_xor_38_nl, loop_DES_rounds_9_xor_38_nl,
      loop_DES_rounds_10_xor_38_nl, loop_DES_rounds_11_xor_38_nl, loop_DES_rounds_12_xor_38_nl,
      loop_DES_rounds_13_xor_38_nl, loop_DES_rounds_14_xor_38_nl, loop_DES_rounds_15_xor_38_nl,
      loop_DES_rounds_16_xor_38_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_49_nl = (reg_input_ftd[4]) ^ (s_output_1_19_16_20_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_6_xor_43_nl = R_23_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign loop_DES_rounds_8_xor_43_nl = R_23_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_9_xor_43_nl = R_23_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_10_xor_43_nl = R_23_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_11_xor_43_nl = R_1_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_12_xor_43_nl = R_23_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_13_xor_43_nl = R_1_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_14_xor_43_nl = R_23_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_15_xor_43_nl = R_1_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_16_xor_43_nl = R_23_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign operator_8_false_1_mux1h_8_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_49_nl,
      loop_DES_rounds_4_xor_97, loop_DES_rounds_5_xor_85, loop_DES_rounds_6_xor_43_nl,
      loop_DES_rounds_2_xor_81, loop_DES_rounds_8_xor_43_nl, loop_DES_rounds_9_xor_43_nl,
      loop_DES_rounds_10_xor_43_nl, loop_DES_rounds_11_xor_43_nl, loop_DES_rounds_12_xor_43_nl,
      loop_DES_rounds_13_xor_43_nl, loop_DES_rounds_14_xor_43_nl, loop_DES_rounds_15_xor_43_nl,
      loop_DES_rounds_16_xor_43_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_50_nl = (key_io_read_key_rsc_cse_63_1_sva[30]) ^ (reg_input_ftd[38])
      ^ (s_output_1_3_0_9_sva[3]);
  assign loop_DES_rounds_4_xor_39_nl = R_27_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_5_xor_39_nl = R_27_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_6_xor_39_nl = R_27_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_7_xor_39_nl = R_27_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_8_xor_39_nl = R_27_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_9_xor_39_nl = R_27_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign loop_DES_rounds_10_xor_39_nl = R_27_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign loop_DES_rounds_11_xor_39_nl = R_27_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_12_xor_39_nl = R_27_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_13_xor_39_nl = R_27_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_14_xor_39_nl = R_27_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_15_xor_39_nl = R_27_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_16_xor_39_nl = R_27_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign operator_8_false_1_mux1h_9_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_50_nl,
      loop_DES_rounds_4_xor_39_nl, loop_DES_rounds_5_xor_39_nl, loop_DES_rounds_6_xor_39_nl,
      loop_DES_rounds_7_xor_39_nl, loop_DES_rounds_8_xor_39_nl, loop_DES_rounds_9_xor_39_nl,
      loop_DES_rounds_10_xor_39_nl, loop_DES_rounds_11_xor_39_nl, loop_DES_rounds_12_xor_39_nl,
      loop_DES_rounds_13_xor_39_nl, loop_DES_rounds_14_xor_39_nl, loop_DES_rounds_15_xor_39_nl,
      loop_DES_rounds_16_xor_39_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_51_nl = (reg_input_ftd[46]) ^ (s_output_1_19_16_50_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_5_xor_40_nl = R_26_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_6_xor_40_nl = R_26_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_7_xor_40_nl = R_26_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_8_xor_40_nl = R_26_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_9_xor_40_nl = R_26_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign loop_DES_rounds_11_xor_40_nl = R_25_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_12_xor_40_nl = R_22_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_13_xor_40_nl = R_25_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_14_xor_40_nl = R_22_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_15_xor_40_nl = R_25_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_16_xor_40_nl = R_22_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign operator_8_false_1_mux1h_10_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_51_nl,
      loop_DES_rounds_4_xor_81, loop_DES_rounds_5_xor_40_nl, loop_DES_rounds_6_xor_40_nl,
      loop_DES_rounds_7_xor_40_nl, loop_DES_rounds_8_xor_40_nl, loop_DES_rounds_9_xor_40_nl,
      loop_DES_rounds_10_xor_81, loop_DES_rounds_11_xor_40_nl, loop_DES_rounds_12_xor_40_nl,
      loop_DES_rounds_13_xor_40_nl, loop_DES_rounds_14_xor_40_nl, loop_DES_rounds_15_xor_40_nl,
      loop_DES_rounds_16_xor_40_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_52_nl = (reg_input_ftd[54]) ^ (s_output_1_3_0_54_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_4_xor_41_nl = R_24_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_5_xor_41_nl = R_22_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_7_xor_41_nl = R_25_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_11_xor_41_nl = R_24_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_14_xor_41_nl = R_15_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_16_xor_41_nl = R_15_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign operator_8_false_1_mux1h_11_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_52_nl,
      loop_DES_rounds_4_xor_41_nl, loop_DES_rounds_5_xor_41_nl, loop_DES_rounds_6_xor_91,
      loop_DES_rounds_7_xor_41_nl, loop_DES_rounds_8_xor_83, loop_DES_rounds_4_xor_81,
      loop_DES_rounds_10_xor_89, loop_DES_rounds_11_xor_41_nl, loop_DES_rounds_9_xor_93,
      loop_DES_rounds_5_xor_83, loop_DES_rounds_14_xor_41_nl, loop_DES_rounds_7_xor_83,
      loop_DES_rounds_16_xor_41_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_53_nl = (key_io_read_key_rsc_cse_63_1_sva[3]) ^ (reg_input_ftd[62])
      ^ (s_output_1_3_0_24_sva[3]);
  assign loop_DES_rounds_4_xor_42_nl = R_24_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_6_xor_42_nl = R_24_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_8_xor_42_nl = R_24_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_9_xor_42_nl = R_24_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_10_xor_42_nl = R_24_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_11_xor_42_nl = R_23_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_12_xor_42_nl = R_24_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_13_xor_42_nl = R_23_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_14_xor_42_nl = R_24_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_15_xor_42_nl = R_23_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign loop_DES_rounds_16_xor_42_nl = R_24_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign operator_8_false_1_mux1h_12_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_53_nl,
      loop_DES_rounds_4_xor_42_nl, loop_DES_rounds_5_xor_83, loop_DES_rounds_6_xor_42_nl,
      loop_DES_rounds_7_xor_83, loop_DES_rounds_8_xor_42_nl, loop_DES_rounds_9_xor_42_nl,
      loop_DES_rounds_10_xor_42_nl, loop_DES_rounds_11_xor_42_nl, loop_DES_rounds_12_xor_42_nl,
      loop_DES_rounds_13_xor_42_nl, loop_DES_rounds_14_xor_42_nl, loop_DES_rounds_15_xor_42_nl,
      loop_DES_rounds_16_xor_42_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign nl_U_ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_10_rg_I_1 = {operator_8_false_1_mux1h_nl
      , operator_8_false_1_mux1h_8_nl , operator_8_false_1_mux1h_9_nl , operator_8_false_1_mux1h_10_nl
      , operator_8_false_1_mux1h_11_nl , operator_8_false_1_mux1h_12_nl};
  wire[0:0] operator_8_false_1_mux1h_1_nl;
  wire[0:0] loop_DES_rounds_1_xor_50_nl;
  wire[0:0] loop_DES_rounds_xor_24_nl;
  wire[0:0] loop_DES_rounds_4_xor_50_nl;
  wire[0:0] loop_DES_rounds_5_xor_50_nl;
  wire[0:0] loop_DES_rounds_7_xor_50_nl;
  wire[0:0] loop_DES_rounds_8_xor_50_nl;
  wire[0:0] loop_DES_rounds_10_xor_50_nl;
  wire[0:0] loop_DES_rounds_12_xor_50_nl;
  wire[0:0] loop_DES_rounds_13_xor_50_nl;
  wire[0:0] loop_DES_rounds_14_xor_50_nl;
  wire[0:0] loop_DES_rounds_15_xor_50_nl;
  wire[0:0] loop_DES_rounds_16_xor_50_nl;
  wire[0:0] operator_8_false_1_mux1h_13_nl;
  wire[0:0] loop_DES_rounds_1_xor_55_nl;
  wire[0:0] loop_DES_rounds_xor_25_nl;
  wire[0:0] loop_DES_rounds_4_xor_55_nl;
  wire[0:0] loop_DES_rounds_5_xor_55_nl;
  wire[0:0] loop_DES_rounds_6_xor_55_nl;
  wire[0:0] loop_DES_rounds_7_xor_55_nl;
  wire[0:0] loop_DES_rounds_8_xor_55_nl;
  wire[0:0] loop_DES_rounds_9_xor_55_nl;
  wire[0:0] loop_DES_rounds_10_xor_55_nl;
  wire[0:0] loop_DES_rounds_11_xor_55_nl;
  wire[0:0] loop_DES_rounds_12_xor_55_nl;
  wire[0:0] loop_DES_rounds_13_xor_55_nl;
  wire[0:0] loop_DES_rounds_14_xor_55_nl;
  wire[0:0] loop_DES_rounds_15_xor_55_nl;
  wire[0:0] operator_8_false_1_mux1h_14_nl;
  wire[0:0] loop_DES_rounds_1_xor_51_nl;
  wire[0:0] loop_DES_rounds_xor_26_nl;
  wire[0:0] loop_DES_rounds_4_xor_51_nl;
  wire[0:0] loop_DES_rounds_5_xor_51_nl;
  wire[0:0] loop_DES_rounds_6_xor_51_nl;
  wire[0:0] loop_DES_rounds_7_xor_51_nl;
  wire[0:0] loop_DES_rounds_8_xor_51_nl;
  wire[0:0] loop_DES_rounds_9_xor_51_nl;
  wire[0:0] loop_DES_rounds_10_xor_51_nl;
  wire[0:0] loop_DES_rounds_11_xor_51_nl;
  wire[0:0] loop_DES_rounds_12_xor_51_nl;
  wire[0:0] loop_DES_rounds_13_xor_51_nl;
  wire[0:0] loop_DES_rounds_14_xor_51_nl;
  wire[0:0] loop_DES_rounds_15_xor_51_nl;
  wire[0:0] loop_DES_rounds_16_xor_51_nl;
  wire[0:0] operator_8_false_1_mux1h_15_nl;
  wire[0:0] loop_DES_rounds_1_xor_52_nl;
  wire[0:0] loop_DES_rounds_xor_27_nl;
  wire[0:0] loop_DES_rounds_4_xor_52_nl;
  wire[0:0] loop_DES_rounds_5_xor_52_nl;
  wire[0:0] loop_DES_rounds_6_xor_52_nl;
  wire[0:0] loop_DES_rounds_7_xor_52_nl;
  wire[0:0] loop_DES_rounds_8_xor_52_nl;
  wire[0:0] loop_DES_rounds_9_xor_52_nl;
  wire[0:0] loop_DES_rounds_10_xor_52_nl;
  wire[0:0] loop_DES_rounds_11_xor_52_nl;
  wire[0:0] loop_DES_rounds_12_xor_52_nl;
  wire[0:0] loop_DES_rounds_13_xor_52_nl;
  wire[0:0] loop_DES_rounds_15_xor_52_nl;
  wire[0:0] loop_DES_rounds_16_xor_52_nl;
  wire[0:0] operator_8_false_1_mux1h_16_nl;
  wire[0:0] loop_DES_rounds_1_xor_53_nl;
  wire[0:0] loop_DES_rounds_xor_28_nl;
  wire[0:0] loop_DES_rounds_4_xor_53_nl;
  wire[0:0] loop_DES_rounds_5_xor_53_nl;
  wire[0:0] loop_DES_rounds_7_xor_53_nl;
  wire[0:0] loop_DES_rounds_8_xor_53_nl;
  wire[0:0] loop_DES_rounds_10_xor_53_nl;
  wire[0:0] loop_DES_rounds_11_xor_53_nl;
  wire[0:0] loop_DES_rounds_12_xor_53_nl;
  wire[0:0] loop_DES_rounds_13_xor_53_nl;
  wire[0:0] loop_DES_rounds_14_xor_53_nl;
  wire[0:0] loop_DES_rounds_15_xor_53_nl;
  wire[0:0] loop_DES_rounds_16_xor_53_nl;
  wire[0:0] operator_8_false_1_mux1h_17_nl;
  wire[0:0] loop_DES_rounds_1_xor_54_nl;
  wire[0:0] loop_DES_rounds_xor_29_nl;
  wire[0:0] loop_DES_rounds_4_xor_54_nl;
  wire[0:0] loop_DES_rounds_5_xor_54_nl;
  wire[0:0] loop_DES_rounds_6_xor_54_nl;
  wire[0:0] loop_DES_rounds_7_xor_54_nl;
  wire[0:0] loop_DES_rounds_8_xor_54_nl;
  wire[0:0] loop_DES_rounds_9_xor_54_nl;
  wire[0:0] loop_DES_rounds_10_xor_54_nl;
  wire[0:0] loop_DES_rounds_11_xor_54_nl;
  wire[0:0] loop_DES_rounds_12_xor_54_nl;
  wire[0:0] loop_DES_rounds_13_xor_54_nl;
  wire[0:0] loop_DES_rounds_14_xor_54_nl;
  wire[0:0] loop_DES_rounds_15_xor_54_nl;
  wire[0:0] loop_DES_rounds_16_xor_54_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_rg_I_1;
  assign loop_DES_rounds_1_xor_50_nl = (input_rsci_idat[29]) ^ (key_rsci_idat[5]);
  assign loop_DES_rounds_xor_24_nl = (key_io_read_key_rsc_cse_63_1_sva[28]) ^ (reg_input_ftd[28])
      ^ (s_output_1_3_0_54_sva[2]);
  assign loop_DES_rounds_4_xor_50_nl = R_20_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_5_xor_50_nl = R_20_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_7_xor_50_nl = R_20_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign loop_DES_rounds_8_xor_50_nl = R_20_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign loop_DES_rounds_10_xor_50_nl = R_20_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_12_xor_50_nl = R_20_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_13_xor_50_nl = R_20_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign loop_DES_rounds_14_xor_50_nl = R_20_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign loop_DES_rounds_15_xor_50_nl = R_20_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign loop_DES_rounds_16_xor_50_nl = R_20_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign operator_8_false_1_mux1h_1_nl = MUX1HOT_s_1_15_2(loop_DES_rounds_1_xor_50_nl,
      loop_DES_rounds_xor_24_nl, loop_DES_rounds_4_xor_50_nl, loop_DES_rounds_5_xor_50_nl,
      loop_DES_rounds_6_xor_87, loop_DES_rounds_7_xor_50_nl, loop_DES_rounds_8_xor_50_nl,
      loop_DES_rounds_9_xor_81, loop_DES_rounds_10_xor_50_nl, loop_DES_rounds_9_xor_89,
      loop_DES_rounds_12_xor_50_nl, loop_DES_rounds_13_xor_50_nl, loop_DES_rounds_14_xor_50_nl,
      loop_DES_rounds_15_xor_50_nl, loop_DES_rounds_16_xor_50_nl, {(fsm_output[0])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9]) , (fsm_output[10]) ,
      (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13]) , (fsm_output[14]) ,
      (fsm_output[15])});
  assign loop_DES_rounds_1_xor_55_nl = (input_rsci_idat[3]) ^ (key_rsci_idat[23]);
  assign loop_DES_rounds_xor_25_nl = (key_io_read_key_rsc_cse_63_1_sva[46]) ^ (reg_input_ftd[2])
      ^ (s_output_1_19_16_20_sva[2]);
  assign loop_DES_rounds_4_xor_55_nl = R_15_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_5_xor_55_nl = R_15_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_6_xor_55_nl = R_15_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_7_xor_55_nl = R_15_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_8_xor_55_nl = R_15_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_9_xor_55_nl = R_15_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign loop_DES_rounds_10_xor_55_nl = R_15_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_11_xor_55_nl = R_15_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_12_xor_55_nl = R_15_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_13_xor_55_nl = R_15_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_14_xor_55_nl = R_15_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_15_xor_55_nl = R_15_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign operator_8_false_1_mux1h_13_nl = MUX1HOT_s_1_15_2(loop_DES_rounds_1_xor_55_nl,
      loop_DES_rounds_xor_25_nl, loop_DES_rounds_4_xor_55_nl, loop_DES_rounds_5_xor_55_nl,
      loop_DES_rounds_6_xor_55_nl, loop_DES_rounds_7_xor_55_nl, loop_DES_rounds_8_xor_55_nl,
      loop_DES_rounds_9_xor_55_nl, loop_DES_rounds_10_xor_55_nl, loop_DES_rounds_11_xor_55_nl,
      loop_DES_rounds_12_xor_55_nl, loop_DES_rounds_13_xor_55_nl, loop_DES_rounds_14_xor_55_nl,
      loop_DES_rounds_15_xor_55_nl, loop_DES_rounds_6_xor_89, {(fsm_output[0]) ,
      (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9]) , (fsm_output[10]) ,
      (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13]) , (fsm_output[14]) ,
      (fsm_output[15])});
  assign loop_DES_rounds_1_xor_51_nl = (input_rsci_idat[37]) ^ (key_rsci_idat[63]);
  assign loop_DES_rounds_xor_26_nl = (key_io_read_key_rsc_cse_63_1_sva[21]) ^ (reg_input_ftd[36])
      ^ (s_output_1_19_16_35_sva[3]);
  assign loop_DES_rounds_4_xor_51_nl = R_19_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign loop_DES_rounds_5_xor_51_nl = R_19_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign loop_DES_rounds_6_xor_51_nl = R_19_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign loop_DES_rounds_7_xor_51_nl = R_19_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_8_xor_51_nl = R_19_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_9_xor_51_nl = R_19_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_10_xor_51_nl = R_19_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_11_xor_51_nl = R_1_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_12_xor_51_nl = R_19_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign loop_DES_rounds_13_xor_51_nl = R_1_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign loop_DES_rounds_14_xor_51_nl = R_19_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign loop_DES_rounds_15_xor_51_nl = R_1_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_16_xor_51_nl = R_19_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign operator_8_false_1_mux1h_14_nl = MUX1HOT_s_1_15_2(loop_DES_rounds_1_xor_51_nl,
      loop_DES_rounds_xor_26_nl, loop_DES_rounds_4_xor_51_nl, loop_DES_rounds_5_xor_51_nl,
      loop_DES_rounds_6_xor_51_nl, loop_DES_rounds_7_xor_51_nl, loop_DES_rounds_8_xor_51_nl,
      loop_DES_rounds_9_xor_51_nl, loop_DES_rounds_10_xor_51_nl, loop_DES_rounds_11_xor_51_nl,
      loop_DES_rounds_12_xor_51_nl, loop_DES_rounds_13_xor_51_nl, loop_DES_rounds_14_xor_51_nl,
      loop_DES_rounds_15_xor_51_nl, loop_DES_rounds_16_xor_51_nl, {(fsm_output[0])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9]) , (fsm_output[10]) ,
      (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13]) , (fsm_output[14]) ,
      (fsm_output[15])});
  assign loop_DES_rounds_1_xor_52_nl = (input_rsci_idat[45]) ^ (key_rsci_idat[28]);
  assign loop_DES_rounds_xor_27_nl = (reg_input_ftd[44]) ^ (s_output_1_3_0_24_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_4_xor_52_nl = R_18_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_5_xor_52_nl = R_27_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_6_xor_52_nl = R_3_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_7_xor_52_nl = R_31_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign loop_DES_rounds_8_xor_52_nl = R_7_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign loop_DES_rounds_9_xor_52_nl = R_27_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_10_xor_52_nl = R_18_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_11_xor_52_nl = R_1_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_12_xor_52_nl = R_3_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign loop_DES_rounds_13_xor_52_nl = R_10_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_15_xor_52_nl = R_31_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_16_xor_52_nl = R_1_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign operator_8_false_1_mux1h_15_nl = MUX1HOT_s_1_15_2(loop_DES_rounds_1_xor_52_nl,
      loop_DES_rounds_xor_27_nl, loop_DES_rounds_4_xor_52_nl, loop_DES_rounds_5_xor_52_nl,
      loop_DES_rounds_6_xor_52_nl, loop_DES_rounds_7_xor_52_nl, loop_DES_rounds_8_xor_52_nl,
      loop_DES_rounds_9_xor_52_nl, loop_DES_rounds_10_xor_52_nl, loop_DES_rounds_11_xor_52_nl,
      loop_DES_rounds_12_xor_52_nl, loop_DES_rounds_13_xor_52_nl, loop_DES_rounds_14_xor_81,
      loop_DES_rounds_15_xor_52_nl, loop_DES_rounds_16_xor_52_nl, {(fsm_output[0])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9]) , (fsm_output[10]) ,
      (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13]) , (fsm_output[14]) ,
      (fsm_output[15])});
  assign loop_DES_rounds_1_xor_53_nl = (input_rsci_idat[53]) ^ (key_rsci_idat[37]);
  assign loop_DES_rounds_xor_28_nl = (reg_input_ftd[52]) ^ (s_output_1_3_0_9_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_4_xor_53_nl = R_15_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_5_xor_53_nl = R_15_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign loop_DES_rounds_7_xor_53_nl = R_15_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign loop_DES_rounds_8_xor_53_nl = R_15_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_10_xor_53_nl = R_15_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_11_xor_53_nl = R_16_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign loop_DES_rounds_12_xor_53_nl = R_16_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign loop_DES_rounds_13_xor_53_nl = R_16_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign loop_DES_rounds_14_xor_53_nl = R_16_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign loop_DES_rounds_15_xor_53_nl = R_16_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_16_xor_53_nl = R_14_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign operator_8_false_1_mux1h_16_nl = MUX1HOT_s_1_15_2(loop_DES_rounds_1_xor_53_nl,
      loop_DES_rounds_xor_28_nl, loop_DES_rounds_4_xor_53_nl, loop_DES_rounds_5_xor_53_nl,
      loop_DES_rounds_6_xor_89, loop_DES_rounds_7_xor_53_nl, loop_DES_rounds_8_xor_53_nl,
      loop_DES_rounds_9_xor_89, loop_DES_rounds_10_xor_53_nl, loop_DES_rounds_11_xor_53_nl,
      loop_DES_rounds_12_xor_53_nl, loop_DES_rounds_13_xor_53_nl, loop_DES_rounds_14_xor_53_nl,
      loop_DES_rounds_15_xor_53_nl, loop_DES_rounds_16_xor_53_nl, {(fsm_output[0])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9]) , (fsm_output[10]) ,
      (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13]) , (fsm_output[14]) ,
      (fsm_output[15])});
  assign loop_DES_rounds_1_xor_54_nl = (input_rsci_idat[61]) ^ (key_rsci_idat[46]);
  assign loop_DES_rounds_xor_29_nl = (key_io_read_key_rsc_cse_63_1_sva[4]) ^ (reg_input_ftd[60])
      ^ (s_output_1_19_16_50_sva[2]);
  assign loop_DES_rounds_4_xor_54_nl = R_16_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_5_xor_54_nl = R_16_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_6_xor_54_nl = R_16_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_7_xor_54_nl = R_16_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_8_xor_54_nl = R_16_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_9_xor_54_nl = R_16_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign loop_DES_rounds_10_xor_54_nl = R_16_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign loop_DES_rounds_11_xor_54_nl = R_15_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign loop_DES_rounds_12_xor_54_nl = R_15_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_13_xor_54_nl = R_15_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_14_xor_54_nl = R_15_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_15_xor_54_nl = R_15_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_16_xor_54_nl = R_15_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign operator_8_false_1_mux1h_17_nl = MUX1HOT_s_1_15_2(loop_DES_rounds_1_xor_54_nl,
      loop_DES_rounds_xor_29_nl, loop_DES_rounds_4_xor_54_nl, loop_DES_rounds_5_xor_54_nl,
      loop_DES_rounds_6_xor_54_nl, loop_DES_rounds_7_xor_54_nl, loop_DES_rounds_8_xor_54_nl,
      loop_DES_rounds_9_xor_54_nl, loop_DES_rounds_10_xor_54_nl, loop_DES_rounds_11_xor_54_nl,
      loop_DES_rounds_12_xor_54_nl, loop_DES_rounds_13_xor_54_nl, loop_DES_rounds_14_xor_54_nl,
      loop_DES_rounds_15_xor_54_nl, loop_DES_rounds_16_xor_54_nl, {(fsm_output[0])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9]) , (fsm_output[10]) ,
      (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13]) , (fsm_output[14]) ,
      (fsm_output[15])});
  assign nl_U_ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_rg_I_1 = {operator_8_false_1_mux1h_1_nl
      , operator_8_false_1_mux1h_13_nl , operator_8_false_1_mux1h_14_nl , operator_8_false_1_mux1h_15_nl
      , operator_8_false_1_mux1h_16_nl , operator_8_false_1_mux1h_17_nl};
  wire[0:0] operator_8_false_1_mux_nl;
  wire[0:0] loop_DES_rounds_2_xor_nl;
  wire[0:0] loop_DES_rounds_16_xor_nl;
  wire[0:0] operator_8_false_1_mux_1_nl;
  wire[0:0] loop_DES_rounds_2_xor_37_nl;
  wire[0:0] loop_DES_rounds_16_xor_37_nl;
  wire[0:0] operator_8_false_1_mux_2_nl;
  wire[0:0] loop_DES_rounds_xor_16_nl;
  wire[0:0] loop_DES_rounds_16_xor_33_nl;
  wire[0:0] operator_8_false_1_mux_3_nl;
  wire[0:0] loop_DES_rounds_xor_17_nl;
  wire[0:0] loop_DES_rounds_16_xor_34_nl;
  wire[0:0] operator_8_false_1_mux_4_nl;
  wire[0:0] operator_8_false_1_mux_5_nl;
  wire[0:0] loop_DES_rounds_2_xor_36_nl;
  wire[0:0] loop_DES_rounds_16_xor_36_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_ce1b43b29576509b87f48de0e64c68b52f_1_rg_I_1;
  assign loop_DES_rounds_2_xor_nl = R_0_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_16_xor_nl = R_0_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign operator_8_false_1_mux_nl = MUX_s_1_2_2(loop_DES_rounds_2_xor_nl, loop_DES_rounds_16_xor_nl,
      fsm_output[15]);
  assign loop_DES_rounds_2_xor_37_nl = R_31_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_16_xor_37_nl = R_27_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign operator_8_false_1_mux_1_nl = MUX_s_1_2_2(loop_DES_rounds_2_xor_37_nl, loop_DES_rounds_16_xor_37_nl,
      fsm_output[15]);
  assign loop_DES_rounds_xor_16_nl = (reg_input_ftd[5]) ^ (s_output_1_19_16_20_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_16_xor_33_nl = R_31_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign operator_8_false_1_mux_2_nl = MUX_s_1_2_2(loop_DES_rounds_xor_16_nl, loop_DES_rounds_16_xor_33_nl,
      fsm_output[15]);
  assign loop_DES_rounds_xor_17_nl = (reg_input_ftd[13]) ^ (ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_17[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign loop_DES_rounds_16_xor_34_nl = R_26_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign operator_8_false_1_mux_3_nl = MUX_s_1_2_2(loop_DES_rounds_xor_17_nl, loop_DES_rounds_16_xor_34_nl,
      fsm_output[15]);
  assign operator_8_false_1_mux_4_nl = MUX_s_1_2_2(loop_DES_rounds_2_xor_89, loop_DES_rounds_14_xor_81,
      fsm_output[15]);
  assign loop_DES_rounds_2_xor_36_nl = R_27_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_16_xor_36_nl = R_28_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign operator_8_false_1_mux_5_nl = MUX_s_1_2_2(loop_DES_rounds_2_xor_36_nl, loop_DES_rounds_16_xor_36_nl,
      fsm_output[15]);
  assign nl_U_ROM_1i6_1o4_ce1b43b29576509b87f48de0e64c68b52f_1_rg_I_1 = {operator_8_false_1_mux_nl
      , operator_8_false_1_mux_1_nl , operator_8_false_1_mux_2_nl , operator_8_false_1_mux_3_nl
      , operator_8_false_1_mux_4_nl , operator_8_false_1_mux_5_nl};
  wire[0:0] operator_8_false_1_mux1h_2_nl;
  wire[0:0] loop_DES_rounds_1_xor_nl;
  wire[0:0] loop_DES_rounds_xor_60_nl;
  wire[0:0] loop_DES_rounds_4_xor_nl;
  wire[0:0] loop_DES_rounds_5_xor_nl;
  wire[0:0] loop_DES_rounds_6_xor_nl;
  wire[0:0] loop_DES_rounds_7_xor_nl;
  wire[0:0] loop_DES_rounds_8_xor_nl;
  wire[0:0] loop_DES_rounds_9_xor_nl;
  wire[0:0] loop_DES_rounds_10_xor_nl;
  wire[0:0] loop_DES_rounds_11_xor_nl;
  wire[0:0] loop_DES_rounds_12_xor_nl;
  wire[0:0] loop_DES_rounds_13_xor_nl;
  wire[0:0] loop_DES_rounds_14_xor_nl;
  wire[0:0] loop_DES_rounds_15_xor_nl;
  wire[0:0] operator_8_false_1_mux1h_18_nl;
  wire[0:0] loop_DES_rounds_1_xor_37_nl;
  wire[0:0] loop_DES_rounds_xor_61_nl;
  wire[0:0] loop_DES_rounds_4_xor_37_nl;
  wire[0:0] loop_DES_rounds_5_xor_37_nl;
  wire[0:0] loop_DES_rounds_6_xor_37_nl;
  wire[0:0] loop_DES_rounds_7_xor_37_nl;
  wire[0:0] loop_DES_rounds_8_xor_37_nl;
  wire[0:0] loop_DES_rounds_10_xor_37_nl;
  wire[0:0] loop_DES_rounds_11_xor_37_nl;
  wire[0:0] loop_DES_rounds_12_xor_37_nl;
  wire[0:0] loop_DES_rounds_13_xor_37_nl;
  wire[0:0] loop_DES_rounds_14_xor_37_nl;
  wire[0:0] loop_DES_rounds_15_xor_37_nl;
  wire[0:0] operator_8_false_1_mux1h_19_nl;
  wire[0:0] loop_DES_rounds_1_xor_33_nl;
  wire[0:0] loop_DES_rounds_xor_62_nl;
  wire[0:0] loop_DES_rounds_4_xor_33_nl;
  wire[0:0] loop_DES_rounds_5_xor_33_nl;
  wire[0:0] loop_DES_rounds_6_xor_33_nl;
  wire[0:0] loop_DES_rounds_7_xor_33_nl;
  wire[0:0] loop_DES_rounds_8_xor_33_nl;
  wire[0:0] loop_DES_rounds_9_xor_33_nl;
  wire[0:0] loop_DES_rounds_10_xor_33_nl;
  wire[0:0] loop_DES_rounds_11_xor_33_nl;
  wire[0:0] loop_DES_rounds_12_xor_33_nl;
  wire[0:0] loop_DES_rounds_13_xor_33_nl;
  wire[0:0] loop_DES_rounds_14_xor_33_nl;
  wire[0:0] loop_DES_rounds_15_xor_33_nl;
  wire[0:0] operator_8_false_1_mux1h_20_nl;
  wire[0:0] loop_DES_rounds_1_xor_34_nl;
  wire[0:0] loop_DES_rounds_xor_63_nl;
  wire[0:0] loop_DES_rounds_4_xor_34_nl;
  wire[0:0] loop_DES_rounds_5_xor_34_nl;
  wire[0:0] loop_DES_rounds_6_xor_34_nl;
  wire[0:0] loop_DES_rounds_7_xor_34_nl;
  wire[0:0] loop_DES_rounds_8_xor_34_nl;
  wire[0:0] loop_DES_rounds_9_xor_34_nl;
  wire[0:0] loop_DES_rounds_10_xor_34_nl;
  wire[0:0] loop_DES_rounds_11_xor_34_nl;
  wire[0:0] loop_DES_rounds_13_xor_34_nl;
  wire[0:0] loop_DES_rounds_14_xor_34_nl;
  wire[0:0] loop_DES_rounds_15_xor_34_nl;
  wire[0:0] operator_8_false_1_mux1h_21_nl;
  wire[0:0] loop_DES_rounds_1_xor_35_nl;
  wire[0:0] loop_DES_rounds_xor_64_nl;
  wire[0:0] loop_DES_rounds_4_xor_35_nl;
  wire[0:0] loop_DES_rounds_5_xor_35_nl;
  wire[0:0] loop_DES_rounds_6_xor_35_nl;
  wire[0:0] loop_DES_rounds_7_xor_35_nl;
  wire[0:0] loop_DES_rounds_8_xor_35_nl;
  wire[0:0] loop_DES_rounds_9_xor_35_nl;
  wire[0:0] loop_DES_rounds_10_xor_35_nl;
  wire[0:0] loop_DES_rounds_12_xor_35_nl;
  wire[0:0] loop_DES_rounds_13_xor_35_nl;
  wire[0:0] loop_DES_rounds_14_xor_35_nl;
  wire[0:0] loop_DES_rounds_15_xor_35_nl;
  wire[0:0] operator_8_false_1_mux1h_22_nl;
  wire[0:0] loop_DES_rounds_1_xor_36_nl;
  wire[0:0] loop_DES_rounds_xor_65_nl;
  wire[0:0] loop_DES_rounds_4_xor_36_nl;
  wire[0:0] loop_DES_rounds_5_xor_36_nl;
  wire[0:0] loop_DES_rounds_6_xor_36_nl;
  wire[0:0] loop_DES_rounds_7_xor_36_nl;
  wire[0:0] loop_DES_rounds_8_xor_36_nl;
  wire[0:0] loop_DES_rounds_9_xor_36_nl;
  wire[0:0] loop_DES_rounds_10_xor_36_nl;
  wire[0:0] loop_DES_rounds_12_xor_36_nl;
  wire[0:0] loop_DES_rounds_13_xor_36_nl;
  wire[0:0] loop_DES_rounds_15_xor_36_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_ce1b43b29576509b87f48de0e64c68b52f_rg_I_1;
  assign loop_DES_rounds_1_xor_nl = (input_rsci_idat[57]) ^ (key_rsci_idat[54]);
  assign loop_DES_rounds_xor_60_nl = (key_io_read_key_rsc_cse_63_1_sva[12]) ^ (reg_input_ftd[56])
      ^ (s_output_1_3_0_54_sva[3]);
  assign loop_DES_rounds_4_xor_nl = R_0_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign loop_DES_rounds_5_xor_nl = R_0_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_6_xor_nl = R_0_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_7_xor_nl = R_0_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_8_xor_nl = R_0_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign loop_DES_rounds_9_xor_nl = R_0_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_10_xor_nl = R_0_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_11_xor_nl = R_0_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_12_xor_nl = R_0_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_13_xor_nl = R_0_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_14_xor_nl = R_0_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign loop_DES_rounds_15_xor_nl = R_0_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign operator_8_false_1_mux1h_2_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_1_xor_nl,
      loop_DES_rounds_xor_60_nl, loop_DES_rounds_4_xor_nl, loop_DES_rounds_5_xor_nl,
      loop_DES_rounds_6_xor_nl, loop_DES_rounds_7_xor_nl, loop_DES_rounds_8_xor_nl,
      loop_DES_rounds_9_xor_nl, loop_DES_rounds_10_xor_nl, loop_DES_rounds_11_xor_nl,
      loop_DES_rounds_12_xor_nl, loop_DES_rounds_13_xor_nl, loop_DES_rounds_14_xor_nl,
      loop_DES_rounds_15_xor_nl, {(fsm_output[0]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])
      , (fsm_output[9]) , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12])
      , (fsm_output[13]) , (fsm_output[14])});
  assign loop_DES_rounds_1_xor_37_nl = (input_rsci_idat[39]) ^ (key_rsci_idat[47]);
  assign loop_DES_rounds_xor_61_nl = (reg_input_ftd[38]) ^ (s_output_1_3_0_9_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_4_xor_37_nl = R_27_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign loop_DES_rounds_5_xor_37_nl = R_27_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign loop_DES_rounds_6_xor_37_nl = R_27_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign loop_DES_rounds_7_xor_37_nl = R_27_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign loop_DES_rounds_8_xor_37_nl = R_27_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_10_xor_37_nl = R_27_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_11_xor_37_nl = R_27_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_12_xor_37_nl = R_27_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_13_xor_37_nl = R_27_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign loop_DES_rounds_14_xor_37_nl = R_27_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign loop_DES_rounds_15_xor_37_nl = R_27_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign operator_8_false_1_mux1h_18_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_1_xor_37_nl,
      loop_DES_rounds_xor_61_nl, loop_DES_rounds_4_xor_37_nl, loop_DES_rounds_5_xor_37_nl,
      loop_DES_rounds_6_xor_37_nl, loop_DES_rounds_7_xor_37_nl, loop_DES_rounds_8_xor_37_nl,
      loop_DES_rounds_9_xor_83, loop_DES_rounds_10_xor_37_nl, loop_DES_rounds_11_xor_37_nl,
      loop_DES_rounds_12_xor_37_nl, loop_DES_rounds_13_xor_37_nl, loop_DES_rounds_14_xor_37_nl,
      loop_DES_rounds_15_xor_37_nl, {(fsm_output[0]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])
      , (fsm_output[9]) , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12])
      , (fsm_output[13]) , (fsm_output[14])});
  assign loop_DES_rounds_1_xor_33_nl = (input_rsci_idat[7]) ^ (key_rsci_idat[13]);
  assign loop_DES_rounds_xor_62_nl = (key_io_read_key_rsc_cse_63_1_sva[36]) ^ (reg_input_ftd[6])
      ^ (s_output_1_19_16_5_sva[0]);
  assign loop_DES_rounds_4_xor_33_nl = R_31_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_5_xor_33_nl = R_31_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_6_xor_33_nl = R_31_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_7_xor_33_nl = R_31_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_8_xor_33_nl = R_31_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_9_xor_33_nl = R_31_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign loop_DES_rounds_10_xor_33_nl = R_31_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_11_xor_33_nl = R_31_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_12_xor_33_nl = R_31_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_13_xor_33_nl = R_31_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_14_xor_33_nl = R_31_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_15_xor_33_nl = R_31_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign operator_8_false_1_mux1h_19_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_1_xor_33_nl,
      loop_DES_rounds_xor_62_nl, loop_DES_rounds_4_xor_33_nl, loop_DES_rounds_5_xor_33_nl,
      loop_DES_rounds_6_xor_33_nl, loop_DES_rounds_7_xor_33_nl, loop_DES_rounds_8_xor_33_nl,
      loop_DES_rounds_9_xor_33_nl, loop_DES_rounds_10_xor_33_nl, loop_DES_rounds_11_xor_33_nl,
      loop_DES_rounds_12_xor_33_nl, loop_DES_rounds_13_xor_33_nl, loop_DES_rounds_14_xor_33_nl,
      loop_DES_rounds_15_xor_33_nl, {(fsm_output[0]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])
      , (fsm_output[9]) , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12])
      , (fsm_output[13]) , (fsm_output[14])});
  assign loop_DES_rounds_1_xor_34_nl = (input_rsci_idat[15]) ^ (key_rsci_idat[30]);
  assign loop_DES_rounds_xor_63_nl = (reg_input_ftd[14]) ^ (s_output_1_19_16_35_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign loop_DES_rounds_4_xor_34_nl = R_3_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign loop_DES_rounds_5_xor_34_nl = R_30_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_6_xor_34_nl = R_3_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_7_xor_34_nl = R_30_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_8_xor_34_nl = R_3_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_9_xor_34_nl = R_30_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_10_xor_34_nl = R_3_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign loop_DES_rounds_11_xor_34_nl = R_3_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign loop_DES_rounds_13_xor_34_nl = R_3_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_14_xor_34_nl = R_26_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_15_xor_34_nl = R_3_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign operator_8_false_1_mux1h_20_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_1_xor_34_nl,
      loop_DES_rounds_xor_63_nl, loop_DES_rounds_4_xor_34_nl, loop_DES_rounds_5_xor_34_nl,
      loop_DES_rounds_6_xor_34_nl, loop_DES_rounds_7_xor_34_nl, loop_DES_rounds_8_xor_34_nl,
      loop_DES_rounds_9_xor_34_nl, loop_DES_rounds_10_xor_34_nl, loop_DES_rounds_11_xor_34_nl,
      loop_DES_rounds_10_xor_81, loop_DES_rounds_13_xor_34_nl, loop_DES_rounds_14_xor_34_nl,
      loop_DES_rounds_15_xor_34_nl, {(fsm_output[0]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])
      , (fsm_output[9]) , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12])
      , (fsm_output[13]) , (fsm_output[14])});
  assign loop_DES_rounds_1_xor_35_nl = (input_rsci_idat[23]) ^ (key_rsci_idat[4]);
  assign loop_DES_rounds_xor_64_nl = (reg_input_ftd[22]) ^ (s_output_1_3_0_24_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign loop_DES_rounds_4_xor_35_nl = R_26_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign loop_DES_rounds_5_xor_35_nl = R_29_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign loop_DES_rounds_6_xor_35_nl = R_29_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_7_xor_35_nl = R_29_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_8_xor_35_nl = R_29_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_9_xor_35_nl = R_29_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign loop_DES_rounds_10_xor_35_nl = R_29_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign loop_DES_rounds_12_xor_35_nl = R_26_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign loop_DES_rounds_13_xor_35_nl = R_28_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_14_xor_35_nl = R_26_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_15_xor_35_nl = R_28_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign operator_8_false_1_mux1h_21_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_1_xor_35_nl,
      loop_DES_rounds_xor_64_nl, loop_DES_rounds_4_xor_35_nl, loop_DES_rounds_5_xor_35_nl,
      loop_DES_rounds_6_xor_35_nl, loop_DES_rounds_7_xor_35_nl, loop_DES_rounds_8_xor_35_nl,
      loop_DES_rounds_9_xor_35_nl, loop_DES_rounds_10_xor_35_nl, loop_DES_rounds_7_xor_85,
      loop_DES_rounds_12_xor_35_nl, loop_DES_rounds_13_xor_35_nl, loop_DES_rounds_14_xor_35_nl,
      loop_DES_rounds_15_xor_35_nl, {(fsm_output[0]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])
      , (fsm_output[9]) , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12])
      , (fsm_output[13]) , (fsm_output[14])});
  assign loop_DES_rounds_1_xor_36_nl = (input_rsci_idat[31]) ^ (key_rsci_idat[15]);
  assign loop_DES_rounds_xor_65_nl = (key_io_read_key_rsc_cse_63_1_sva[38]) ^ (reg_input_ftd[30])
      ^ (s_output_1_3_0_39_sva[3]);
  assign loop_DES_rounds_4_xor_36_nl = R_28_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_5_xor_36_nl = R_28_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_6_xor_36_nl = R_28_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign loop_DES_rounds_7_xor_36_nl = R_28_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign loop_DES_rounds_8_xor_36_nl = R_28_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign loop_DES_rounds_9_xor_36_nl = R_28_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_10_xor_36_nl = R_28_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_12_xor_36_nl = R_28_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_13_xor_36_nl = R_27_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_15_xor_36_nl = R_27_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[27]);
  assign operator_8_false_1_mux1h_22_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_1_xor_36_nl,
      loop_DES_rounds_xor_65_nl, loop_DES_rounds_4_xor_36_nl, loop_DES_rounds_5_xor_36_nl,
      loop_DES_rounds_6_xor_36_nl, loop_DES_rounds_7_xor_36_nl, loop_DES_rounds_8_xor_36_nl,
      loop_DES_rounds_9_xor_36_nl, loop_DES_rounds_10_xor_36_nl, loop_DES_rounds_9_xor_83,
      loop_DES_rounds_12_xor_36_nl, loop_DES_rounds_13_xor_36_nl, loop_DES_rounds_2_xor_89,
      loop_DES_rounds_15_xor_36_nl, {(fsm_output[0]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])
      , (fsm_output[9]) , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12])
      , (fsm_output[13]) , (fsm_output[14])});
  assign nl_U_ROM_1i6_1o4_ce1b43b29576509b87f48de0e64c68b52f_rg_I_1 = {operator_8_false_1_mux1h_2_nl
      , operator_8_false_1_mux1h_18_nl , operator_8_false_1_mux1h_19_nl , operator_8_false_1_mux1h_20_nl
      , operator_8_false_1_mux1h_21_nl , operator_8_false_1_mux1h_22_nl};
  wire[0:0] operator_8_false_1_mux1h_3_nl;
  wire[0:0] loop_DES_rounds_xor_30_nl;
  wire[0:0] loop_DES_rounds_5_xor_68_nl;
  wire[0:0] loop_DES_rounds_6_xor_68_nl;
  wire[0:0] loop_DES_rounds_7_xor_68_nl;
  wire[0:0] loop_DES_rounds_8_xor_68_nl;
  wire[0:0] loop_DES_rounds_9_xor_68_nl;
  wire[0:0] loop_DES_rounds_10_xor_68_nl;
  wire[0:0] loop_DES_rounds_13_xor_68_nl;
  wire[0:0] loop_DES_rounds_14_xor_68_nl;
  wire[0:0] loop_DES_rounds_15_xor_68_nl;
  wire[0:0] loop_DES_rounds_16_xor_68_nl;
  wire[0:0] operator_8_false_1_mux1h_23_nl;
  wire[0:0] loop_DES_rounds_xor_31_nl;
  wire[0:0] loop_DES_rounds_5_xor_73_nl;
  wire[0:0] loop_DES_rounds_6_xor_73_nl;
  wire[0:0] loop_DES_rounds_7_xor_73_nl;
  wire[0:0] loop_DES_rounds_8_xor_73_nl;
  wire[0:0] loop_DES_rounds_9_xor_73_nl;
  wire[0:0] loop_DES_rounds_10_xor_73_nl;
  wire[0:0] loop_DES_rounds_12_xor_73_nl;
  wire[0:0] loop_DES_rounds_13_xor_73_nl;
  wire[0:0] loop_DES_rounds_14_xor_73_nl;
  wire[0:0] loop_DES_rounds_16_xor_73_nl;
  wire[0:0] operator_8_false_1_mux1h_24_nl;
  wire[0:0] loop_DES_rounds_xor_32_nl;
  wire[0:0] loop_DES_rounds_4_xor_69_nl;
  wire[0:0] loop_DES_rounds_5_xor_69_nl;
  wire[0:0] loop_DES_rounds_6_xor_69_nl;
  wire[0:0] loop_DES_rounds_7_xor_69_nl;
  wire[0:0] loop_DES_rounds_9_xor_69_nl;
  wire[0:0] loop_DES_rounds_10_xor_69_nl;
  wire[0:0] loop_DES_rounds_11_xor_69_nl;
  wire[0:0] loop_DES_rounds_12_xor_69_nl;
  wire[0:0] loop_DES_rounds_13_xor_69_nl;
  wire[0:0] loop_DES_rounds_14_xor_69_nl;
  wire[0:0] loop_DES_rounds_15_xor_69_nl;
  wire[0:0] loop_DES_rounds_16_xor_69_nl;
  wire[0:0] operator_8_false_1_mux1h_25_nl;
  wire[0:0] loop_DES_rounds_xor_33_nl;
  wire[0:0] loop_DES_rounds_5_xor_70_nl;
  wire[0:0] loop_DES_rounds_6_xor_70_nl;
  wire[0:0] loop_DES_rounds_7_xor_70_nl;
  wire[0:0] loop_DES_rounds_8_xor_70_nl;
  wire[0:0] loop_DES_rounds_9_xor_70_nl;
  wire[0:0] loop_DES_rounds_10_xor_70_nl;
  wire[0:0] loop_DES_rounds_11_xor_70_nl;
  wire[0:0] loop_DES_rounds_12_xor_70_nl;
  wire[0:0] loop_DES_rounds_13_xor_70_nl;
  wire[0:0] loop_DES_rounds_14_xor_70_nl;
  wire[0:0] loop_DES_rounds_15_xor_70_nl;
  wire[0:0] loop_DES_rounds_16_xor_70_nl;
  wire[0:0] operator_8_false_1_mux1h_26_nl;
  wire[0:0] loop_DES_rounds_xor_34_nl;
  wire[0:0] loop_DES_rounds_5_xor_71_nl;
  wire[0:0] loop_DES_rounds_6_xor_71_nl;
  wire[0:0] loop_DES_rounds_7_xor_71_nl;
  wire[0:0] loop_DES_rounds_8_xor_71_nl;
  wire[0:0] loop_DES_rounds_9_xor_71_nl;
  wire[0:0] loop_DES_rounds_10_xor_71_nl;
  wire[0:0] loop_DES_rounds_11_xor_71_nl;
  wire[0:0] loop_DES_rounds_12_xor_71_nl;
  wire[0:0] loop_DES_rounds_13_xor_71_nl;
  wire[0:0] loop_DES_rounds_14_xor_71_nl;
  wire[0:0] loop_DES_rounds_15_xor_71_nl;
  wire[0:0] loop_DES_rounds_16_xor_71_nl;
  wire[0:0] operator_8_false_1_mux1h_27_nl;
  wire[0:0] loop_DES_rounds_xor_35_nl;
  wire[0:0] loop_DES_rounds_4_xor_72_nl;
  wire[0:0] loop_DES_rounds_5_xor_72_nl;
  wire[0:0] loop_DES_rounds_6_xor_72_nl;
  wire[0:0] loop_DES_rounds_7_xor_72_nl;
  wire[0:0] loop_DES_rounds_8_xor_72_nl;
  wire[0:0] loop_DES_rounds_9_xor_72_nl;
  wire[0:0] loop_DES_rounds_10_xor_72_nl;
  wire[0:0] loop_DES_rounds_11_xor_72_nl;
  wire[0:0] loop_DES_rounds_12_xor_72_nl;
  wire[0:0] loop_DES_rounds_13_xor_72_nl;
  wire[0:0] loop_DES_rounds_14_xor_72_nl;
  wire[0:0] loop_DES_rounds_15_xor_72_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_10_rg_I_1;
  assign loop_DES_rounds_xor_30_nl = (reg_input_ftd[58]) ^ (s_output_1_19_16_50_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_5_xor_68_nl = R_8_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_6_xor_68_nl = R_7_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_7_xor_68_nl = R_8_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_8_xor_68_nl = R_7_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_9_xor_68_nl = R_8_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_10_xor_68_nl = R_7_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_13_xor_68_nl = R_7_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_14_xor_68_nl = R_7_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_15_xor_68_nl = R_7_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_16_xor_68_nl = R_7_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign operator_8_false_1_mux1h_3_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_30_nl,
      loop_DES_rounds_4_xor_85, loop_DES_rounds_5_xor_68_nl, loop_DES_rounds_6_xor_68_nl,
      loop_DES_rounds_7_xor_68_nl, loop_DES_rounds_8_xor_68_nl, loop_DES_rounds_9_xor_68_nl,
      loop_DES_rounds_10_xor_68_nl, loop_DES_rounds_9_xor_87, loop_DES_rounds_10_xor_87,
      loop_DES_rounds_13_xor_68_nl, loop_DES_rounds_14_xor_68_nl, loop_DES_rounds_15_xor_68_nl,
      loop_DES_rounds_16_xor_68_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_31_nl = (key_io_read_key_rsc_cse_63_1_sva[0]) ^ (reg_input_ftd[32])
      ^ (s_output_1_3_0_39_sva[2]);
  assign loop_DES_rounds_5_xor_73_nl = R_3_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_6_xor_73_nl = R_3_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_7_xor_73_nl = R_3_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_8_xor_73_nl = R_3_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_9_xor_73_nl = R_3_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign loop_DES_rounds_10_xor_73_nl = R_3_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_12_xor_73_nl = R_3_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_13_xor_73_nl = R_3_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_14_xor_73_nl = R_3_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_16_xor_73_nl = R_3_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign operator_8_false_1_mux1h_23_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_31_nl,
      loop_DES_rounds_4_xor_95, loop_DES_rounds_5_xor_73_nl, loop_DES_rounds_6_xor_73_nl,
      loop_DES_rounds_7_xor_73_nl, loop_DES_rounds_8_xor_73_nl, loop_DES_rounds_9_xor_73_nl,
      loop_DES_rounds_10_xor_73_nl, loop_DES_rounds_2_xor_91, loop_DES_rounds_12_xor_73_nl,
      loop_DES_rounds_13_xor_73_nl, loop_DES_rounds_14_xor_73_nl, loop_DES_rounds_9_xor_91,
      loop_DES_rounds_16_xor_73_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_32_nl = (key_io_read_key_rsc_cse_63_1_sva[35]) ^ (reg_input_ftd[0])
      ^ (s_output_1_3_0_24_sva[1]);
  assign loop_DES_rounds_4_xor_69_nl = R_7_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_5_xor_69_nl = R_7_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_6_xor_69_nl = R_7_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_7_xor_69_nl = R_7_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_9_xor_69_nl = R_7_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign loop_DES_rounds_10_xor_69_nl = R_7_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_11_xor_69_nl = R_7_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign loop_DES_rounds_12_xor_69_nl = R_7_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_13_xor_69_nl = R_7_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_14_xor_69_nl = R_7_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_15_xor_69_nl = R_7_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_16_xor_69_nl = R_7_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign operator_8_false_1_mux1h_24_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_32_nl,
      loop_DES_rounds_4_xor_69_nl, loop_DES_rounds_5_xor_69_nl, loop_DES_rounds_6_xor_69_nl,
      loop_DES_rounds_7_xor_69_nl, loop_DES_rounds_2_xor_85, loop_DES_rounds_9_xor_69_nl,
      loop_DES_rounds_10_xor_69_nl, loop_DES_rounds_11_xor_69_nl, loop_DES_rounds_12_xor_69_nl,
      loop_DES_rounds_13_xor_69_nl, loop_DES_rounds_14_xor_69_nl, loop_DES_rounds_15_xor_69_nl,
      loop_DES_rounds_16_xor_69_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_33_nl = (reg_input_ftd[8]) ^ (s_output_1_19_16_5_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_5_xor_70_nl = R_1_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_6_xor_70_nl = R_6_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_7_xor_70_nl = R_1_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_8_xor_70_nl = R_6_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_9_xor_70_nl = R_1_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_10_xor_70_nl = R_6_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_11_xor_70_nl = R_30_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_12_xor_70_nl = R_29_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_13_xor_70_nl = R_30_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_14_xor_70_nl = R_29_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign loop_DES_rounds_15_xor_70_nl = R_30_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_16_xor_70_nl = R_29_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign operator_8_false_1_mux1h_25_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_33_nl,
      loop_DES_rounds_4_xor_89, loop_DES_rounds_5_xor_70_nl, loop_DES_rounds_6_xor_70_nl,
      loop_DES_rounds_7_xor_70_nl, loop_DES_rounds_8_xor_70_nl, loop_DES_rounds_9_xor_70_nl,
      loop_DES_rounds_10_xor_70_nl, loop_DES_rounds_11_xor_70_nl, loop_DES_rounds_12_xor_70_nl,
      loop_DES_rounds_13_xor_70_nl, loop_DES_rounds_14_xor_70_nl, loop_DES_rounds_15_xor_70_nl,
      loop_DES_rounds_16_xor_70_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_34_nl = (reg_input_ftd[16]) ^ (s_output_1_3_0_9_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_5_xor_71_nl = R_0_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign loop_DES_rounds_6_xor_71_nl = R_4_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_7_xor_71_nl = R_0_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign loop_DES_rounds_8_xor_71_nl = R_4_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_9_xor_71_nl = R_0_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_10_xor_71_nl = R_4_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_11_xor_71_nl = R_4_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_12_xor_71_nl = R_29_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_13_xor_71_nl = R_4_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_14_xor_71_nl = R_29_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_15_xor_71_nl = R_4_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_16_xor_71_nl = R_26_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign operator_8_false_1_mux1h_26_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_34_nl,
      loop_DES_rounds_4_xor_83, loop_DES_rounds_5_xor_71_nl, loop_DES_rounds_6_xor_71_nl,
      loop_DES_rounds_7_xor_71_nl, loop_DES_rounds_8_xor_71_nl, loop_DES_rounds_9_xor_71_nl,
      loop_DES_rounds_10_xor_71_nl, loop_DES_rounds_11_xor_71_nl, loop_DES_rounds_12_xor_71_nl,
      loop_DES_rounds_13_xor_71_nl, loop_DES_rounds_14_xor_71_nl, loop_DES_rounds_15_xor_71_nl,
      loop_DES_rounds_16_xor_71_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_35_nl = (key_io_read_key_rsc_cse_63_1_sva[9]) ^ (reg_input_ftd[24])
      ^ (s_output_1_19_16_35_sva[2]);
  assign loop_DES_rounds_4_xor_72_nl = R_31_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign loop_DES_rounds_5_xor_72_nl = R_4_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_6_xor_72_nl = R_31_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_7_xor_72_nl = R_4_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_8_xor_72_nl = R_31_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_9_xor_72_nl = R_4_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_10_xor_72_nl = R_31_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_11_xor_72_nl = R_31_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_12_xor_72_nl = R_4_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_13_xor_72_nl = R_31_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_14_xor_72_nl = R_4_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_15_xor_72_nl = R_31_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign operator_8_false_1_mux1h_27_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_35_nl,
      loop_DES_rounds_4_xor_72_nl, loop_DES_rounds_5_xor_72_nl, loop_DES_rounds_6_xor_72_nl,
      loop_DES_rounds_7_xor_72_nl, loop_DES_rounds_8_xor_72_nl, loop_DES_rounds_9_xor_72_nl,
      loop_DES_rounds_10_xor_72_nl, loop_DES_rounds_11_xor_72_nl, loop_DES_rounds_12_xor_72_nl,
      loop_DES_rounds_13_xor_72_nl, loop_DES_rounds_14_xor_72_nl, loop_DES_rounds_15_xor_72_nl,
      loop_DES_rounds_4_xor_83, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign nl_U_ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_10_rg_I_1 = {operator_8_false_1_mux1h_3_nl
      , operator_8_false_1_mux1h_23_nl , operator_8_false_1_mux1h_24_nl , operator_8_false_1_mux1h_25_nl
      , operator_8_false_1_mux1h_26_nl , operator_8_false_1_mux1h_27_nl};
  wire[0:0] operator_8_false_1_mux1h_4_nl;
  wire[0:0] loop_DES_rounds_xor_54_nl;
  wire[0:0] loop_DES_rounds_4_xor_56_nl;
  wire[0:0] loop_DES_rounds_5_xor_56_nl;
  wire[0:0] loop_DES_rounds_6_xor_56_nl;
  wire[0:0] loop_DES_rounds_7_xor_56_nl;
  wire[0:0] loop_DES_rounds_8_xor_56_nl;
  wire[0:0] loop_DES_rounds_9_xor_56_nl;
  wire[0:0] loop_DES_rounds_10_xor_56_nl;
  wire[0:0] loop_DES_rounds_12_xor_56_nl;
  wire[0:0] loop_DES_rounds_14_xor_56_nl;
  wire[0:0] loop_DES_rounds_15_xor_56_nl;
  wire[0:0] operator_8_false_1_mux1h_28_nl;
  wire[0:0] loop_DES_rounds_xor_55_nl;
  wire[0:0] loop_DES_rounds_4_xor_61_nl;
  wire[0:0] loop_DES_rounds_5_xor_61_nl;
  wire[0:0] loop_DES_rounds_7_xor_61_nl;
  wire[0:0] loop_DES_rounds_8_xor_61_nl;
  wire[0:0] loop_DES_rounds_10_xor_61_nl;
  wire[0:0] loop_DES_rounds_11_xor_61_nl;
  wire[0:0] loop_DES_rounds_12_xor_61_nl;
  wire[0:0] loop_DES_rounds_13_xor_61_nl;
  wire[0:0] loop_DES_rounds_14_xor_61_nl;
  wire[0:0] loop_DES_rounds_15_xor_61_nl;
  wire[0:0] loop_DES_rounds_16_xor_61_nl;
  wire[0:0] operator_8_false_1_mux1h_29_nl;
  wire[0:0] loop_DES_rounds_xor_56_nl;
  wire[0:0] loop_DES_rounds_4_xor_57_nl;
  wire[0:0] loop_DES_rounds_6_xor_57_nl;
  wire[0:0] loop_DES_rounds_8_xor_57_nl;
  wire[0:0] loop_DES_rounds_9_xor_57_nl;
  wire[0:0] loop_DES_rounds_12_xor_57_nl;
  wire[0:0] loop_DES_rounds_13_xor_57_nl;
  wire[0:0] loop_DES_rounds_14_xor_57_nl;
  wire[0:0] loop_DES_rounds_15_xor_57_nl;
  wire[0:0] loop_DES_rounds_16_xor_57_nl;
  wire[0:0] operator_8_false_1_mux1h_30_nl;
  wire[0:0] loop_DES_rounds_xor_57_nl;
  wire[0:0] loop_DES_rounds_4_xor_58_nl;
  wire[0:0] loop_DES_rounds_5_xor_58_nl;
  wire[0:0] loop_DES_rounds_6_xor_58_nl;
  wire[0:0] loop_DES_rounds_7_xor_58_nl;
  wire[0:0] loop_DES_rounds_8_xor_58_nl;
  wire[0:0] loop_DES_rounds_9_xor_58_nl;
  wire[0:0] loop_DES_rounds_10_xor_58_nl;
  wire[0:0] loop_DES_rounds_11_xor_58_nl;
  wire[0:0] loop_DES_rounds_12_xor_58_nl;
  wire[0:0] loop_DES_rounds_13_xor_58_nl;
  wire[0:0] loop_DES_rounds_14_xor_58_nl;
  wire[0:0] loop_DES_rounds_15_xor_58_nl;
  wire[0:0] operator_8_false_1_mux1h_31_nl;
  wire[0:0] loop_DES_rounds_xor_58_nl;
  wire[0:0] loop_DES_rounds_4_xor_59_nl;
  wire[0:0] loop_DES_rounds_5_xor_59_nl;
  wire[0:0] loop_DES_rounds_7_xor_59_nl;
  wire[0:0] loop_DES_rounds_11_xor_59_nl;
  wire[0:0] loop_DES_rounds_12_xor_59_nl;
  wire[0:0] loop_DES_rounds_13_xor_59_nl;
  wire[0:0] loop_DES_rounds_14_xor_59_nl;
  wire[0:0] loop_DES_rounds_15_xor_59_nl;
  wire[0:0] operator_8_false_1_mux1h_32_nl;
  wire[0:0] loop_DES_rounds_xor_59_nl;
  wire[0:0] loop_DES_rounds_4_xor_60_nl;
  wire[0:0] loop_DES_rounds_5_xor_60_nl;
  wire[0:0] loop_DES_rounds_6_xor_60_nl;
  wire[0:0] loop_DES_rounds_7_xor_60_nl;
  wire[0:0] loop_DES_rounds_9_xor_60_nl;
  wire[0:0] loop_DES_rounds_11_xor_60_nl;
  wire[0:0] loop_DES_rounds_12_xor_60_nl;
  wire[0:0] loop_DES_rounds_14_xor_60_nl;
  wire[0:0] loop_DES_rounds_15_xor_60_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_10_rg_I_1;
  assign loop_DES_rounds_xor_54_nl = (key_io_read_key_rsc_cse_63_1_sva[2]) ^ (reg_input_ftd[60])
      ^ (s_output_1_19_16_50_sva[2]);
  assign loop_DES_rounds_4_xor_56_nl = R_16_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_5_xor_56_nl = R_16_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_6_xor_56_nl = R_16_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_7_xor_56_nl = R_16_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_8_xor_56_nl = R_16_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_9_xor_56_nl = R_16_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_10_xor_56_nl = R_16_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_12_xor_56_nl = R_15_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_14_xor_56_nl = R_15_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_15_xor_56_nl = R_15_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign operator_8_false_1_mux1h_4_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_54_nl,
      loop_DES_rounds_4_xor_56_nl, loop_DES_rounds_5_xor_56_nl, loop_DES_rounds_6_xor_56_nl,
      loop_DES_rounds_7_xor_56_nl, loop_DES_rounds_8_xor_56_nl, loop_DES_rounds_9_xor_56_nl,
      loop_DES_rounds_10_xor_56_nl, loop_DES_rounds_5_xor_81, loop_DES_rounds_12_xor_56_nl,
      loop_DES_rounds_7_xor_87, loop_DES_rounds_14_xor_56_nl, loop_DES_rounds_15_xor_56_nl,
      loop_DES_rounds_10_xor_83, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_55_nl = (key_io_read_key_rsc_cse_63_1_sva[16]) ^ (reg_input_ftd[34])
      ^ (s_output_1_3_0_9_sva[0]);
  assign loop_DES_rounds_4_xor_61_nl = R_11_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_5_xor_61_nl = R_11_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_7_xor_61_nl = R_11_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_8_xor_61_nl = R_11_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_10_xor_61_nl = R_11_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_11_xor_61_nl = R_11_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_12_xor_61_nl = R_11_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_13_xor_61_nl = R_11_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_14_xor_61_nl = R_11_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_15_xor_61_nl = R_11_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_16_xor_61_nl = R_11_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign operator_8_false_1_mux1h_28_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_55_nl,
      loop_DES_rounds_4_xor_61_nl, loop_DES_rounds_5_xor_61_nl, loop_DES_rounds_6_xor_83,
      loop_DES_rounds_7_xor_61_nl, loop_DES_rounds_8_xor_61_nl, loop_DES_rounds_9_xor_85,
      loop_DES_rounds_10_xor_61_nl, loop_DES_rounds_11_xor_61_nl, loop_DES_rounds_12_xor_61_nl,
      loop_DES_rounds_13_xor_61_nl, loop_DES_rounds_14_xor_61_nl, loop_DES_rounds_15_xor_61_nl,
      loop_DES_rounds_16_xor_61_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_56_nl = (key_io_read_key_rsc_cse_63_1_sva[59]) ^ (reg_input_ftd[2])
      ^ (s_output_1_19_16_20_sva[2]);
  assign loop_DES_rounds_4_xor_57_nl = R_15_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_6_xor_57_nl = R_15_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_8_xor_57_nl = R_15_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_9_xor_57_nl = R_15_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_12_xor_57_nl = R_15_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_13_xor_57_nl = R_15_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_14_xor_57_nl = R_15_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_15_xor_57_nl = R_15_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_16_xor_57_nl = R_15_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign operator_8_false_1_mux1h_29_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_56_nl,
      loop_DES_rounds_4_xor_57_nl, loop_DES_rounds_5_xor_81, loop_DES_rounds_6_xor_57_nl,
      loop_DES_rounds_7_xor_87, loop_DES_rounds_8_xor_57_nl, loop_DES_rounds_9_xor_57_nl,
      loop_DES_rounds_10_xor_83, loop_DES_rounds_2_xor_87, loop_DES_rounds_12_xor_57_nl,
      loop_DES_rounds_13_xor_57_nl, loop_DES_rounds_14_xor_57_nl, loop_DES_rounds_15_xor_57_nl,
      loop_DES_rounds_16_xor_57_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_57_nl = (reg_input_ftd[10]) ^ (s_output_1_19_16_35_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_4_xor_58_nl = R_14_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_5_xor_58_nl = R_31_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_6_xor_58_nl = R_7_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_7_xor_58_nl = R_1_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_8_xor_58_nl = R_10_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_9_xor_58_nl = R_1_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_10_xor_58_nl = R_12_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_11_xor_58_nl = R_1_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_12_xor_58_nl = R_31_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_13_xor_58_nl = R_1_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_14_xor_58_nl = R_1_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_15_xor_58_nl = R_10_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign operator_8_false_1_mux1h_30_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_57_nl,
      loop_DES_rounds_4_xor_58_nl, loop_DES_rounds_5_xor_58_nl, loop_DES_rounds_6_xor_58_nl,
      loop_DES_rounds_7_xor_58_nl, loop_DES_rounds_8_xor_58_nl, loop_DES_rounds_9_xor_58_nl,
      loop_DES_rounds_10_xor_58_nl, loop_DES_rounds_11_xor_58_nl, loop_DES_rounds_12_xor_58_nl,
      loop_DES_rounds_13_xor_58_nl, loop_DES_rounds_14_xor_58_nl, loop_DES_rounds_15_xor_58_nl,
      loop_DES_rounds_2_xor_93, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_58_nl = (reg_input_ftd[18]) ^ (s_output_1_3_0_39_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_4_xor_59_nl = R_12_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_5_xor_59_nl = R_20_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_7_xor_59_nl = R_27_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_11_xor_59_nl = R_12_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_12_xor_59_nl = R_24_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_13_xor_59_nl = R_12_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_14_xor_59_nl = R_3_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_15_xor_59_nl = R_12_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign operator_8_false_1_mux1h_31_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_58_nl,
      loop_DES_rounds_4_xor_59_nl, loop_DES_rounds_5_xor_59_nl, loop_DES_rounds_6_xor_93,
      loop_DES_rounds_7_xor_59_nl, loop_DES_rounds_8_xor_89, loop_DES_rounds_9_xor_91,
      loop_DES_rounds_10_xor_85, loop_DES_rounds_11_xor_59_nl, loop_DES_rounds_12_xor_59_nl,
      loop_DES_rounds_13_xor_59_nl, loop_DES_rounds_14_xor_59_nl, loop_DES_rounds_15_xor_59_nl,
      loop_DES_rounds_6_xor_83, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_59_nl = (key_io_read_key_rsc_cse_63_1_sva[50]) ^ (reg_input_ftd[26])
      ^ (s_output_1_19_16_5_sva[2]);
  assign loop_DES_rounds_4_xor_60_nl = R_11_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_5_xor_60_nl = R_12_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_6_xor_60_nl = R_11_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_7_xor_60_nl = R_12_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_9_xor_60_nl = R_12_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_11_xor_60_nl = R_11_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_12_xor_60_nl = R_12_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign loop_DES_rounds_14_xor_60_nl = R_12_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_15_xor_60_nl = R_11_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign operator_8_false_1_mux1h_32_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_59_nl,
      loop_DES_rounds_4_xor_60_nl, loop_DES_rounds_5_xor_60_nl, loop_DES_rounds_6_xor_60_nl,
      loop_DES_rounds_7_xor_60_nl, loop_DES_rounds_8_xor_85, loop_DES_rounds_9_xor_60_nl,
      loop_DES_rounds_4_xor_91, loop_DES_rounds_11_xor_60_nl, loop_DES_rounds_12_xor_60_nl,
      loop_DES_rounds_9_xor_85, loop_DES_rounds_14_xor_60_nl, loop_DES_rounds_15_xor_60_nl,
      loop_DES_rounds_6_xor_93, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign nl_U_ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_10_rg_I_1 = {operator_8_false_1_mux1h_4_nl
      , operator_8_false_1_mux1h_28_nl , operator_8_false_1_mux1h_29_nl , operator_8_false_1_mux1h_30_nl
      , operator_8_false_1_mux1h_31_nl , operator_8_false_1_mux1h_32_nl};
  wire[0:0] operator_8_false_1_mux1h_5_nl;
  wire[0:0] loop_DES_rounds_xor_36_nl;
  wire[0:0] loop_DES_rounds_4_xor_44_nl;
  wire[0:0] loop_DES_rounds_5_xor_44_nl;
  wire[0:0] loop_DES_rounds_6_xor_44_nl;
  wire[0:0] loop_DES_rounds_7_xor_44_nl;
  wire[0:0] loop_DES_rounds_8_xor_44_nl;
  wire[0:0] loop_DES_rounds_9_xor_44_nl;
  wire[0:0] loop_DES_rounds_10_xor_44_nl;
  wire[0:0] loop_DES_rounds_11_xor_44_nl;
  wire[0:0] operator_8_false_1_mux1h_33_nl;
  wire[0:0] loop_DES_rounds_xor_37_nl;
  wire[0:0] loop_DES_rounds_4_xor_49_nl;
  wire[0:0] loop_DES_rounds_5_xor_49_nl;
  wire[0:0] loop_DES_rounds_6_xor_49_nl;
  wire[0:0] loop_DES_rounds_7_xor_49_nl;
  wire[0:0] loop_DES_rounds_8_xor_49_nl;
  wire[0:0] loop_DES_rounds_9_xor_49_nl;
  wire[0:0] loop_DES_rounds_10_xor_49_nl;
  wire[0:0] loop_DES_rounds_11_xor_49_nl;
  wire[0:0] loop_DES_rounds_12_xor_49_nl;
  wire[0:0] loop_DES_rounds_13_xor_49_nl;
  wire[0:0] loop_DES_rounds_14_xor_49_nl;
  wire[0:0] loop_DES_rounds_15_xor_49_nl;
  wire[0:0] loop_DES_rounds_16_xor_49_nl;
  wire[0:0] operator_8_false_1_mux1h_34_nl;
  wire[0:0] loop_DES_rounds_xor_38_nl;
  wire[0:0] loop_DES_rounds_5_xor_45_nl;
  wire[0:0] loop_DES_rounds_6_xor_45_nl;
  wire[0:0] loop_DES_rounds_7_xor_45_nl;
  wire[0:0] loop_DES_rounds_8_xor_45_nl;
  wire[0:0] loop_DES_rounds_9_xor_45_nl;
  wire[0:0] loop_DES_rounds_10_xor_45_nl;
  wire[0:0] loop_DES_rounds_11_xor_45_nl;
  wire[0:0] loop_DES_rounds_12_xor_45_nl;
  wire[0:0] loop_DES_rounds_13_xor_45_nl;
  wire[0:0] loop_DES_rounds_15_xor_45_nl;
  wire[0:0] loop_DES_rounds_16_xor_45_nl;
  wire[0:0] operator_8_false_1_mux1h_35_nl;
  wire[0:0] loop_DES_rounds_xor_39_nl;
  wire[0:0] loop_DES_rounds_5_xor_46_nl;
  wire[0:0] loop_DES_rounds_6_xor_46_nl;
  wire[0:0] loop_DES_rounds_7_xor_46_nl;
  wire[0:0] loop_DES_rounds_8_xor_46_nl;
  wire[0:0] loop_DES_rounds_10_xor_46_nl;
  wire[0:0] loop_DES_rounds_11_xor_46_nl;
  wire[0:0] loop_DES_rounds_12_xor_46_nl;
  wire[0:0] loop_DES_rounds_13_xor_46_nl;
  wire[0:0] loop_DES_rounds_14_xor_46_nl;
  wire[0:0] loop_DES_rounds_15_xor_46_nl;
  wire[0:0] loop_DES_rounds_16_xor_46_nl;
  wire[0:0] operator_8_false_1_mux1h_36_nl;
  wire[0:0] loop_DES_rounds_xor_40_nl;
  wire[0:0] loop_DES_rounds_4_xor_47_nl;
  wire[0:0] loop_DES_rounds_5_xor_47_nl;
  wire[0:0] loop_DES_rounds_6_xor_47_nl;
  wire[0:0] loop_DES_rounds_7_xor_47_nl;
  wire[0:0] loop_DES_rounds_9_xor_47_nl;
  wire[0:0] loop_DES_rounds_10_xor_47_nl;
  wire[0:0] loop_DES_rounds_11_xor_47_nl;
  wire[0:0] loop_DES_rounds_12_xor_47_nl;
  wire[0:0] loop_DES_rounds_13_xor_47_nl;
  wire[0:0] loop_DES_rounds_14_xor_47_nl;
  wire[0:0] loop_DES_rounds_16_xor_47_nl;
  wire[0:0] operator_8_false_1_mux1h_37_nl;
  wire[0:0] loop_DES_rounds_xor_41_nl;
  wire[0:0] loop_DES_rounds_4_xor_48_nl;
  wire[0:0] loop_DES_rounds_5_xor_48_nl;
  wire[0:0] loop_DES_rounds_6_xor_48_nl;
  wire[0:0] loop_DES_rounds_7_xor_48_nl;
  wire[0:0] loop_DES_rounds_8_xor_48_nl;
  wire[0:0] loop_DES_rounds_9_xor_48_nl;
  wire[0:0] loop_DES_rounds_10_xor_48_nl;
  wire[0:0] loop_DES_rounds_11_xor_48_nl;
  wire[0:0] loop_DES_rounds_12_xor_48_nl;
  wire[0:0] loop_DES_rounds_13_xor_48_nl;
  wire[0:0] loop_DES_rounds_14_xor_48_nl;
  wire[0:0] loop_DES_rounds_15_xor_48_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_10_rg_I_1;
  assign loop_DES_rounds_xor_36_nl = (key_io_read_key_rsc_cse_63_1_sva[19]) ^ (reg_input_ftd[62])
      ^ (s_output_1_3_0_24_sva[3]);
  assign loop_DES_rounds_4_xor_44_nl = R_24_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_5_xor_44_nl = R_24_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_6_xor_44_nl = R_24_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_7_xor_44_nl = R_24_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_8_xor_44_nl = R_24_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_9_xor_44_nl = R_24_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_10_xor_44_nl = R_24_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_11_xor_44_nl = R_23_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign operator_8_false_1_mux1h_5_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_36_nl,
      loop_DES_rounds_4_xor_44_nl, loop_DES_rounds_5_xor_44_nl, loop_DES_rounds_6_xor_44_nl,
      loop_DES_rounds_7_xor_44_nl, loop_DES_rounds_8_xor_44_nl, loop_DES_rounds_9_xor_44_nl,
      loop_DES_rounds_10_xor_44_nl, loop_DES_rounds_11_xor_44_nl, loop_DES_rounds_6_xor_91,
      loop_DES_rounds_5_xor_85, loop_DES_rounds_8_xor_83, loop_DES_rounds_2_xor_81,
      loop_DES_rounds_10_xor_89, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_37_nl = (key_io_read_key_rsc_cse_63_1_sva[29]) ^ (reg_input_ftd[36])
      ^ (s_output_1_19_16_35_sva[3]);
  assign loop_DES_rounds_4_xor_49_nl = R_19_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_5_xor_49_nl = R_19_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_6_xor_49_nl = R_19_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_7_xor_49_nl = R_19_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign loop_DES_rounds_8_xor_49_nl = R_19_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_9_xor_49_nl = R_19_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_10_xor_49_nl = R_19_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_11_xor_49_nl = R_1_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_12_xor_49_nl = R_19_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_13_xor_49_nl = R_1_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_14_xor_49_nl = R_19_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_15_xor_49_nl = R_1_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_16_xor_49_nl = R_19_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign operator_8_false_1_mux1h_33_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_37_nl,
      loop_DES_rounds_4_xor_49_nl, loop_DES_rounds_5_xor_49_nl, loop_DES_rounds_6_xor_49_nl,
      loop_DES_rounds_7_xor_49_nl, loop_DES_rounds_8_xor_49_nl, loop_DES_rounds_9_xor_49_nl,
      loop_DES_rounds_10_xor_49_nl, loop_DES_rounds_11_xor_49_nl, loop_DES_rounds_12_xor_49_nl,
      loop_DES_rounds_13_xor_49_nl, loop_DES_rounds_14_xor_49_nl, loop_DES_rounds_15_xor_49_nl,
      loop_DES_rounds_16_xor_49_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_38_nl = (key_io_read_key_rsc_cse_63_1_sva[52]) ^ (reg_input_ftd[4])
      ^ (s_output_1_19_16_20_sva[3]);
  assign loop_DES_rounds_5_xor_45_nl = R_23_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_6_xor_45_nl = R_23_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_7_xor_45_nl = R_23_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_8_xor_45_nl = R_23_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_9_xor_45_nl = R_23_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_10_xor_45_nl = R_23_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_11_xor_45_nl = R_1_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_12_xor_45_nl = R_23_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_13_xor_45_nl = R_1_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_15_xor_45_nl = R_1_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_16_xor_45_nl = R_23_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign operator_8_false_1_mux1h_34_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_38_nl,
      loop_DES_rounds_2_xor_83, loop_DES_rounds_5_xor_45_nl, loop_DES_rounds_6_xor_45_nl,
      loop_DES_rounds_7_xor_45_nl, loop_DES_rounds_8_xor_45_nl, loop_DES_rounds_9_xor_45_nl,
      loop_DES_rounds_10_xor_45_nl, loop_DES_rounds_11_xor_45_nl, loop_DES_rounds_12_xor_45_nl,
      loop_DES_rounds_13_xor_45_nl, loop_DES_rounds_4_xor_97, loop_DES_rounds_15_xor_45_nl,
      loop_DES_rounds_16_xor_45_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_39_nl = (reg_input_ftd[12]) ^ (s_output_1_19_16_5_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_5_xor_46_nl = R_11_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign loop_DES_rounds_6_xor_46_nl = R_21_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_7_xor_46_nl = R_15_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_8_xor_46_nl = R_22_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_10_xor_46_nl = R_22_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_11_xor_46_nl = R_10_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_12_xor_46_nl = R_21_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_13_xor_46_nl = R_21_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_14_xor_46_nl = R_21_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[5]);
  assign loop_DES_rounds_15_xor_46_nl = R_21_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[21]);
  assign loop_DES_rounds_16_xor_46_nl = R_21_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign operator_8_false_1_mux1h_35_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_39_nl,
      loop_DES_rounds_4_xor_93, loop_DES_rounds_5_xor_46_nl, loop_DES_rounds_6_xor_46_nl,
      loop_DES_rounds_7_xor_46_nl, loop_DES_rounds_8_xor_46_nl, loop_DES_rounds_9_xor_93,
      loop_DES_rounds_10_xor_46_nl, loop_DES_rounds_11_xor_46_nl, loop_DES_rounds_12_xor_46_nl,
      loop_DES_rounds_13_xor_46_nl, loop_DES_rounds_14_xor_46_nl, loop_DES_rounds_15_xor_46_nl,
      loop_DES_rounds_16_xor_46_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_40_nl = (reg_input_ftd[20]) ^ (s_output_1_3_0_39_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_4_xor_47_nl = R_21_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_5_xor_47_nl = R_1_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_6_xor_47_nl = R_10_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[45]);
  assign loop_DES_rounds_7_xor_47_nl = R_21_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_9_xor_47_nl = R_21_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_10_xor_47_nl = R_21_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_11_xor_47_nl = R_20_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_12_xor_47_nl = R_2_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_13_xor_47_nl = R_20_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  assign loop_DES_rounds_14_xor_47_nl = R_2_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_16_xor_47_nl = R_2_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign operator_8_false_1_mux1h_36_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_40_nl,
      loop_DES_rounds_4_xor_47_nl, loop_DES_rounds_5_xor_47_nl, loop_DES_rounds_6_xor_47_nl,
      loop_DES_rounds_7_xor_47_nl, loop_DES_rounds_4_xor_93, loop_DES_rounds_9_xor_47_nl,
      loop_DES_rounds_10_xor_47_nl, loop_DES_rounds_11_xor_47_nl, loop_DES_rounds_12_xor_47_nl,
      loop_DES_rounds_13_xor_47_nl, loop_DES_rounds_14_xor_47_nl, loop_DES_rounds_9_xor_81,
      loop_DES_rounds_16_xor_47_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_41_nl = (key_io_read_key_rsc_cse_63_1_sva[14]) ^ (reg_input_ftd[28])
      ^ (s_output_1_3_0_54_sva[2]);
  assign loop_DES_rounds_4_xor_48_nl = R_20_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign loop_DES_rounds_5_xor_48_nl = R_20_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[46]);
  assign loop_DES_rounds_6_xor_48_nl = R_20_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[62]);
  assign loop_DES_rounds_7_xor_48_nl = R_20_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[13]);
  assign loop_DES_rounds_8_xor_48_nl = R_20_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[29]);
  assign loop_DES_rounds_9_xor_48_nl = R_20_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[37]);
  assign loop_DES_rounds_10_xor_48_nl = R_20_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign loop_DES_rounds_11_xor_48_nl = R_20_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[4]);
  assign loop_DES_rounds_12_xor_48_nl = R_20_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[20]);
  assign loop_DES_rounds_13_xor_48_nl = R_20_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_14_xor_48_nl = R_20_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_15_xor_48_nl = R_20_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign operator_8_false_1_mux1h_37_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_41_nl,
      loop_DES_rounds_4_xor_48_nl, loop_DES_rounds_5_xor_48_nl, loop_DES_rounds_6_xor_48_nl,
      loop_DES_rounds_7_xor_48_nl, loop_DES_rounds_8_xor_48_nl, loop_DES_rounds_9_xor_48_nl,
      loop_DES_rounds_10_xor_48_nl, loop_DES_rounds_11_xor_48_nl, loop_DES_rounds_12_xor_48_nl,
      loop_DES_rounds_13_xor_48_nl, loop_DES_rounds_14_xor_48_nl, loop_DES_rounds_15_xor_48_nl,
      loop_DES_rounds_6_xor_87, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign nl_U_ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_10_rg_I_1 = {operator_8_false_1_mux1h_5_nl
      , operator_8_false_1_mux1h_33_nl , operator_8_false_1_mux1h_34_nl , operator_8_false_1_mux1h_35_nl
      , operator_8_false_1_mux1h_36_nl , operator_8_false_1_mux1h_37_nl};
  wire[0:0] operator_8_false_1_mux1h_6_nl;
  wire[0:0] loop_DES_rounds_xor_13_nl;
  wire[0:0] loop_DES_rounds_xor_42_nl;
  wire[0:0] loop_DES_rounds_5_xor_62_nl;
  wire[0:0] loop_DES_rounds_7_xor_62_nl;
  wire[0:0] loop_DES_rounds_8_xor_62_nl;
  wire[0:0] loop_DES_rounds_9_xor_62_nl;
  wire[0:0] loop_DES_rounds_10_xor_62_nl;
  wire[0:0] loop_DES_rounds_11_xor_62_nl;
  wire[0:0] loop_DES_rounds_13_xor_62_nl;
  wire[0:0] loop_DES_rounds_14_xor_62_nl;
  wire[0:0] loop_DES_rounds_15_xor_62_nl;
  wire[0:0] loop_DES_rounds_16_xor_62_nl;
  wire[0:0] operator_8_false_1_mux1h_38_nl;
  wire[0:0] loop_DES_rounds_2_xor_67_nl;
  wire[0:0] loop_DES_rounds_xor_43_nl;
  wire[0:0] loop_DES_rounds_8_xor_67_nl;
  wire[0:0] loop_DES_rounds_11_xor_67_nl;
  wire[0:0] loop_DES_rounds_12_xor_67_nl;
  wire[0:0] loop_DES_rounds_13_xor_67_nl;
  wire[0:0] loop_DES_rounds_14_xor_67_nl;
  wire[0:0] loop_DES_rounds_15_xor_67_nl;
  wire[0:0] loop_DES_rounds_16_xor_67_nl;
  wire[0:0] operator_8_false_1_mux1h_39_nl;
  wire[0:0] loop_DES_rounds_2_xor_63_nl;
  wire[0:0] loop_DES_rounds_xor_44_nl;
  wire[0:0] loop_DES_rounds_4_xor_63_nl;
  wire[0:0] loop_DES_rounds_5_xor_63_nl;
  wire[0:0] loop_DES_rounds_6_xor_63_nl;
  wire[0:0] loop_DES_rounds_7_xor_63_nl;
  wire[0:0] loop_DES_rounds_8_xor_63_nl;
  wire[0:0] loop_DES_rounds_9_xor_63_nl;
  wire[0:0] loop_DES_rounds_10_xor_63_nl;
  wire[0:0] loop_DES_rounds_11_xor_63_nl;
  wire[0:0] loop_DES_rounds_13_xor_63_nl;
  wire[0:0] loop_DES_rounds_14_xor_63_nl;
  wire[0:0] loop_DES_rounds_15_xor_63_nl;
  wire[0:0] operator_8_false_1_mux1h_40_nl;
  wire[0:0] loop_DES_rounds_2_xor_64_nl;
  wire[0:0] loop_DES_rounds_xor_45_nl;
  wire[0:0] loop_DES_rounds_4_xor_64_nl;
  wire[0:0] loop_DES_rounds_5_xor_64_nl;
  wire[0:0] loop_DES_rounds_6_xor_64_nl;
  wire[0:0] loop_DES_rounds_7_xor_64_nl;
  wire[0:0] loop_DES_rounds_8_xor_64_nl;
  wire[0:0] loop_DES_rounds_9_xor_64_nl;
  wire[0:0] loop_DES_rounds_10_xor_64_nl;
  wire[0:0] loop_DES_rounds_11_xor_64_nl;
  wire[0:0] loop_DES_rounds_13_xor_64_nl;
  wire[0:0] loop_DES_rounds_14_xor_64_nl;
  wire[0:0] loop_DES_rounds_16_xor_64_nl;
  wire[0:0] operator_8_false_1_mux1h_41_nl;
  wire[0:0] loop_DES_rounds_xor_46_nl;
  wire[0:0] loop_DES_rounds_4_xor_65_nl;
  wire[0:0] loop_DES_rounds_5_xor_65_nl;
  wire[0:0] loop_DES_rounds_6_xor_65_nl;
  wire[0:0] loop_DES_rounds_7_xor_65_nl;
  wire[0:0] loop_DES_rounds_8_xor_65_nl;
  wire[0:0] loop_DES_rounds_9_xor_65_nl;
  wire[0:0] loop_DES_rounds_10_xor_65_nl;
  wire[0:0] loop_DES_rounds_11_xor_65_nl;
  wire[0:0] loop_DES_rounds_12_xor_65_nl;
  wire[0:0] loop_DES_rounds_13_xor_65_nl;
  wire[0:0] loop_DES_rounds_14_xor_65_nl;
  wire[0:0] loop_DES_rounds_15_xor_65_nl;
  wire[0:0] operator_8_false_1_mux1h_42_nl;
  wire[0:0] loop_DES_rounds_xor_47_nl;
  wire[0:0] loop_DES_rounds_4_xor_66_nl;
  wire[0:0] loop_DES_rounds_5_xor_66_nl;
  wire[0:0] loop_DES_rounds_6_xor_66_nl;
  wire[0:0] loop_DES_rounds_7_xor_66_nl;
  wire[0:0] loop_DES_rounds_9_xor_66_nl;
  wire[0:0] loop_DES_rounds_11_xor_66_nl;
  wire[0:0] loop_DES_rounds_16_xor_66_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_1_rg_I_1;
  assign loop_DES_rounds_xor_13_nl = (reg_input_ftd[25]) ^ (s_output_1_19_16_20_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_xor_42_nl = (reg_input_ftd[26]) ^ (s_output_1_19_16_5_sva[2])
      ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_5_xor_62_nl = R_12_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_7_xor_62_nl = R_12_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_8_xor_62_nl = R_11_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_9_xor_62_nl = R_12_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_10_xor_62_nl = R_11_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_11_xor_62_nl = R_11_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_13_xor_62_nl = R_11_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_14_xor_62_nl = R_12_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_15_xor_62_nl = R_11_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_16_xor_62_nl = R_12_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign operator_8_false_1_mux1h_6_nl = MUX1HOT_s_1_15_2(loop_DES_rounds_xor_13_nl,
      loop_DES_rounds_xor_42_nl, loop_DES_rounds_4_xor_91, loop_DES_rounds_5_xor_62_nl,
      loop_DES_rounds_6_xor_81, loop_DES_rounds_7_xor_62_nl, loop_DES_rounds_8_xor_62_nl,
      loop_DES_rounds_9_xor_62_nl, loop_DES_rounds_10_xor_62_nl, loop_DES_rounds_11_xor_62_nl,
      loop_DES_rounds_8_xor_89, loop_DES_rounds_13_xor_62_nl, loop_DES_rounds_14_xor_62_nl,
      loop_DES_rounds_15_xor_62_nl, loop_DES_rounds_16_xor_62_nl, {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9]) , (fsm_output[10]) ,
      (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13]) , (fsm_output[14]) ,
      (fsm_output[15])});
  assign loop_DES_rounds_2_xor_67_nl = R_7_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_xor_43_nl = (key_io_read_key_rsc_cse_63_1_sva[58]) ^ (reg_input_ftd[0])
      ^ (s_output_1_3_0_24_sva[1]);
  assign loop_DES_rounds_8_xor_67_nl = R_7_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_11_xor_67_nl = R_7_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_12_xor_67_nl = R_7_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_13_xor_67_nl = R_7_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_14_xor_67_nl = R_7_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_15_xor_67_nl = R_7_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_16_xor_67_nl = R_7_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign operator_8_false_1_mux1h_38_nl = MUX1HOT_s_1_15_2(loop_DES_rounds_2_xor_67_nl,
      loop_DES_rounds_xor_43_nl, loop_DES_rounds_4_xor_87, loop_DES_rounds_5_xor_89,
      loop_DES_rounds_6_xor_85, loop_DES_rounds_7_xor_81, loop_DES_rounds_8_xor_67_nl,
      loop_DES_rounds_9_xor_87, loop_DES_rounds_10_xor_87, loop_DES_rounds_11_xor_67_nl,
      loop_DES_rounds_12_xor_67_nl, loop_DES_rounds_13_xor_67_nl, loop_DES_rounds_14_xor_67_nl,
      loop_DES_rounds_15_xor_67_nl, loop_DES_rounds_16_xor_67_nl, {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9]) , (fsm_output[10]) ,
      (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13]) , (fsm_output[14]) ,
      (fsm_output[15])});
  assign loop_DES_rounds_2_xor_63_nl = R_11_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_xor_44_nl = (key_io_read_key_rsc_cse_63_1_sva[57]) ^ (reg_input_ftd[34])
      ^ (s_output_1_3_0_9_sva[0]);
  assign loop_DES_rounds_4_xor_63_nl = R_11_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_5_xor_63_nl = R_11_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_6_xor_63_nl = R_11_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_7_xor_63_nl = R_11_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_8_xor_63_nl = R_11_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_9_xor_63_nl = R_11_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_10_xor_63_nl = R_11_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_11_xor_63_nl = R_11_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_13_xor_63_nl = R_11_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_14_xor_63_nl = R_11_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_15_xor_63_nl = R_11_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign operator_8_false_1_mux1h_39_nl = MUX1HOT_s_1_15_2(loop_DES_rounds_2_xor_63_nl,
      loop_DES_rounds_xor_44_nl, loop_DES_rounds_4_xor_63_nl, loop_DES_rounds_5_xor_63_nl,
      loop_DES_rounds_6_xor_63_nl, loop_DES_rounds_7_xor_63_nl, loop_DES_rounds_8_xor_63_nl,
      loop_DES_rounds_9_xor_63_nl, loop_DES_rounds_10_xor_63_nl, loop_DES_rounds_11_xor_63_nl,
      loop_DES_rounds_8_xor_85, loop_DES_rounds_13_xor_63_nl, loop_DES_rounds_14_xor_63_nl,
      loop_DES_rounds_15_xor_63_nl, loop_DES_rounds_6_xor_81, {(fsm_output[1]) ,
      (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9]) , (fsm_output[10]) ,
      (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13]) , (fsm_output[14]) ,
      (fsm_output[15])});
  assign loop_DES_rounds_2_xor_64_nl = R_10_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_xor_45_nl = (reg_input_ftd[42]) ^ (s_output_1_3_0_54_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_4_xor_64_nl = R_10_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_5_xor_64_nl = R_1_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_6_xor_64_nl = R_1_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_7_xor_64_nl = R_1_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_8_xor_64_nl = R_0_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_9_xor_64_nl = R_10_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_10_xor_64_nl = R_1_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign loop_DES_rounds_11_xor_64_nl = R_10_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_13_xor_64_nl = R_1_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_14_xor_64_nl = R_1_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_16_xor_64_nl = R_0_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign operator_8_false_1_mux1h_40_nl = MUX1HOT_s_1_15_2(loop_DES_rounds_2_xor_64_nl,
      loop_DES_rounds_xor_45_nl, loop_DES_rounds_4_xor_64_nl, loop_DES_rounds_5_xor_64_nl,
      loop_DES_rounds_6_xor_64_nl, loop_DES_rounds_7_xor_64_nl, loop_DES_rounds_8_xor_64_nl,
      loop_DES_rounds_9_xor_64_nl, loop_DES_rounds_10_xor_64_nl, loop_DES_rounds_11_xor_64_nl,
      loop_DES_rounds_5_xor_87, loop_DES_rounds_13_xor_64_nl, loop_DES_rounds_14_xor_64_nl,
      loop_DES_rounds_8_xor_87, loop_DES_rounds_16_xor_64_nl, {(fsm_output[1]) ,
      (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9]) , (fsm_output[10]) ,
      (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13]) , (fsm_output[14]) ,
      (fsm_output[15])});
  assign loop_DES_rounds_xor_46_nl = (reg_input_ftd[50]) ^ (s_output_1_19_16_20_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_4_xor_65_nl = R_6_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_5_xor_65_nl = R_9_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_6_xor_65_nl = R_14_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_7_xor_65_nl = R_9_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_8_xor_65_nl = R_14_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_9_xor_65_nl = R_9_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_10_xor_65_nl = R_14_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_11_xor_65_nl = R_8_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign loop_DES_rounds_12_xor_65_nl = R_0_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_13_xor_65_nl = R_8_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign loop_DES_rounds_14_xor_65_nl = R_0_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_15_xor_65_nl = R_8_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign operator_8_false_1_mux1h_41_nl = MUX1HOT_s_1_15_2(loop_DES_rounds_2_xor_95,
      loop_DES_rounds_xor_46_nl, loop_DES_rounds_4_xor_65_nl, loop_DES_rounds_5_xor_65_nl,
      loop_DES_rounds_6_xor_65_nl, loop_DES_rounds_7_xor_65_nl, loop_DES_rounds_8_xor_65_nl,
      loop_DES_rounds_9_xor_65_nl, loop_DES_rounds_10_xor_65_nl, loop_DES_rounds_11_xor_65_nl,
      loop_DES_rounds_12_xor_65_nl, loop_DES_rounds_13_xor_65_nl, loop_DES_rounds_14_xor_65_nl,
      loop_DES_rounds_15_xor_65_nl, loop_DES_rounds_4_xor_89, {(fsm_output[1]) ,
      (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9]) , (fsm_output[10]) ,
      (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13]) , (fsm_output[14]) ,
      (fsm_output[15])});
  assign loop_DES_rounds_xor_47_nl = (key_io_read_key_rsc_cse_63_1_sva[1]) ^ (reg_input_ftd[58])
      ^ (s_output_1_19_16_50_sva[3]);
  assign loop_DES_rounds_4_xor_66_nl = R_7_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_5_xor_66_nl = R_8_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_6_xor_66_nl = R_7_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_7_xor_66_nl = R_8_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_9_xor_66_nl = R_8_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_11_xor_66_nl = R_7_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_16_xor_66_nl = R_7_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign operator_8_false_1_mux1h_42_nl = MUX1HOT_s_1_15_2(loop_DES_rounds_2_xor_85,
      loop_DES_rounds_xor_47_nl, loop_DES_rounds_4_xor_66_nl, loop_DES_rounds_5_xor_66_nl,
      loop_DES_rounds_6_xor_66_nl, loop_DES_rounds_7_xor_66_nl, loop_DES_rounds_2_xor_95,
      loop_DES_rounds_9_xor_66_nl, loop_DES_rounds_4_xor_85, loop_DES_rounds_11_xor_66_nl,
      loop_DES_rounds_4_xor_87, loop_DES_rounds_5_xor_89, loop_DES_rounds_6_xor_85,
      loop_DES_rounds_7_xor_81, loop_DES_rounds_16_xor_66_nl, {(fsm_output[1]) ,
      (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9]) , (fsm_output[10]) ,
      (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13]) , (fsm_output[14]) ,
      (fsm_output[15])});
  assign nl_U_ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_1_rg_I_1 = {operator_8_false_1_mux1h_6_nl
      , operator_8_false_1_mux1h_38_nl , operator_8_false_1_mux1h_39_nl , operator_8_false_1_mux1h_40_nl
      , operator_8_false_1_mux1h_41_nl , operator_8_false_1_mux1h_42_nl};
  wire[0:0] operator_8_false_1_mux1h_7_nl;
  wire[0:0] loop_DES_rounds_xor_18_nl;
  wire[0:0] loop_DES_rounds_4_xor_74_nl;
  wire[0:0] loop_DES_rounds_5_xor_74_nl;
  wire[0:0] loop_DES_rounds_6_xor_74_nl;
  wire[0:0] loop_DES_rounds_7_xor_74_nl;
  wire[0:0] loop_DES_rounds_9_xor_74_nl;
  wire[0:0] loop_DES_rounds_10_xor_74_nl;
  wire[0:0] loop_DES_rounds_11_xor_74_nl;
  wire[0:0] loop_DES_rounds_12_xor_74_nl;
  wire[0:0] loop_DES_rounds_13_xor_74_nl;
  wire[0:0] loop_DES_rounds_14_xor_74_nl;
  wire[0:0] loop_DES_rounds_15_xor_74_nl;
  wire[0:0] loop_DES_rounds_16_xor_74_nl;
  wire[0:0] operator_8_false_1_mux1h_43_nl;
  wire[0:0] loop_DES_rounds_xor_19_nl;
  wire[0:0] loop_DES_rounds_4_xor_79_nl;
  wire[0:0] loop_DES_rounds_5_xor_79_nl;
  wire[0:0] loop_DES_rounds_6_xor_79_nl;
  wire[0:0] loop_DES_rounds_7_xor_79_nl;
  wire[0:0] loop_DES_rounds_8_xor_79_nl;
  wire[0:0] loop_DES_rounds_9_xor_79_nl;
  wire[0:0] loop_DES_rounds_10_xor_79_nl;
  wire[0:0] loop_DES_rounds_11_xor_79_nl;
  wire[0:0] loop_DES_rounds_12_xor_79_nl;
  wire[0:0] loop_DES_rounds_13_xor_79_nl;
  wire[0:0] loop_DES_rounds_14_xor_79_nl;
  wire[0:0] loop_DES_rounds_15_xor_79_nl;
  wire[0:0] operator_8_false_1_mux1h_44_nl;
  wire[0:0] loop_DES_rounds_xor_20_nl;
  wire[0:0] loop_DES_rounds_4_xor_75_nl;
  wire[0:0] loop_DES_rounds_5_xor_75_nl;
  wire[0:0] loop_DES_rounds_6_xor_75_nl;
  wire[0:0] loop_DES_rounds_7_xor_75_nl;
  wire[0:0] loop_DES_rounds_8_xor_75_nl;
  wire[0:0] loop_DES_rounds_9_xor_75_nl;
  wire[0:0] loop_DES_rounds_11_xor_75_nl;
  wire[0:0] loop_DES_rounds_12_xor_75_nl;
  wire[0:0] loop_DES_rounds_13_xor_75_nl;
  wire[0:0] loop_DES_rounds_14_xor_75_nl;
  wire[0:0] loop_DES_rounds_15_xor_75_nl;
  wire[0:0] loop_DES_rounds_16_xor_75_nl;
  wire[0:0] operator_8_false_1_mux1h_45_nl;
  wire[0:0] loop_DES_rounds_xor_21_nl;
  wire[0:0] loop_DES_rounds_4_xor_76_nl;
  wire[0:0] loop_DES_rounds_5_xor_76_nl;
  wire[0:0] loop_DES_rounds_6_xor_76_nl;
  wire[0:0] loop_DES_rounds_7_xor_76_nl;
  wire[0:0] loop_DES_rounds_8_xor_76_nl;
  wire[0:0] loop_DES_rounds_9_xor_76_nl;
  wire[0:0] loop_DES_rounds_10_xor_76_nl;
  wire[0:0] loop_DES_rounds_11_xor_76_nl;
  wire[0:0] loop_DES_rounds_12_xor_76_nl;
  wire[0:0] loop_DES_rounds_13_xor_76_nl;
  wire[0:0] loop_DES_rounds_14_xor_76_nl;
  wire[0:0] loop_DES_rounds_15_xor_76_nl;
  wire[0:0] loop_DES_rounds_16_xor_76_nl;
  wire[0:0] operator_8_false_1_mux1h_46_nl;
  wire[0:0] loop_DES_rounds_xor_22_nl;
  wire[0:0] loop_DES_rounds_4_xor_77_nl;
  wire[0:0] loop_DES_rounds_6_xor_77_nl;
  wire[0:0] loop_DES_rounds_7_xor_77_nl;
  wire[0:0] loop_DES_rounds_9_xor_77_nl;
  wire[0:0] loop_DES_rounds_10_xor_77_nl;
  wire[0:0] loop_DES_rounds_11_xor_77_nl;
  wire[0:0] loop_DES_rounds_12_xor_77_nl;
  wire[0:0] loop_DES_rounds_13_xor_77_nl;
  wire[0:0] loop_DES_rounds_14_xor_77_nl;
  wire[0:0] loop_DES_rounds_15_xor_77_nl;
  wire[0:0] loop_DES_rounds_16_xor_77_nl;
  wire[0:0] operator_8_false_1_mux1h_47_nl;
  wire[0:0] loop_DES_rounds_xor_23_nl;
  wire[0:0] loop_DES_rounds_4_xor_78_nl;
  wire[0:0] loop_DES_rounds_5_xor_78_nl;
  wire[0:0] loop_DES_rounds_6_xor_78_nl;
  wire[0:0] loop_DES_rounds_7_xor_78_nl;
  wire[0:0] loop_DES_rounds_8_xor_78_nl;
  wire[0:0] loop_DES_rounds_9_xor_78_nl;
  wire[0:0] loop_DES_rounds_10_xor_78_nl;
  wire[0:0] loop_DES_rounds_11_xor_78_nl;
  wire[0:0] loop_DES_rounds_12_xor_78_nl;
  wire[0:0] loop_DES_rounds_13_xor_78_nl;
  wire[0:0] loop_DES_rounds_15_xor_78_nl;
  wire[0:0] loop_DES_rounds_16_xor_78_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_10_rg_I_1;
  assign loop_DES_rounds_xor_18_nl = (key_io_read_key_rsc_cse_63_1_sva[42]) ^ (reg_input_ftd[24])
      ^ (s_output_1_19_16_35_sva[2]);
  assign loop_DES_rounds_4_xor_74_nl = R_31_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_5_xor_74_nl = R_4_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_6_xor_74_nl = R_31_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_7_xor_74_nl = R_4_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_9_xor_74_nl = R_4_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_10_xor_74_nl = R_31_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_11_xor_74_nl = R_31_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_12_xor_74_nl = R_4_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_13_xor_74_nl = R_31_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_14_xor_74_nl = R_4_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_15_xor_74_nl = R_31_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_16_xor_74_nl = R_4_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign operator_8_false_1_mux1h_7_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_18_nl,
      loop_DES_rounds_4_xor_74_nl, loop_DES_rounds_5_xor_74_nl, loop_DES_rounds_6_xor_74_nl,
      loop_DES_rounds_7_xor_74_nl, loop_DES_rounds_8_xor_81, loop_DES_rounds_9_xor_74_nl,
      loop_DES_rounds_10_xor_74_nl, loop_DES_rounds_11_xor_74_nl, loop_DES_rounds_12_xor_74_nl,
      loop_DES_rounds_13_xor_74_nl, loop_DES_rounds_14_xor_74_nl, loop_DES_rounds_15_xor_74_nl,
      loop_DES_rounds_16_xor_74_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_19_nl = (reg_input_ftd[6]) ^ (s_output_1_19_16_5_sva[0])
      ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign loop_DES_rounds_4_xor_79_nl = R_31_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[9]);
  assign loop_DES_rounds_5_xor_79_nl = R_31_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign loop_DES_rounds_6_xor_79_nl = R_31_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_7_xor_79_nl = R_31_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_8_xor_79_nl = R_31_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_9_xor_79_nl = R_31_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_10_xor_79_nl = R_31_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_11_xor_79_nl = R_31_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_12_xor_79_nl = R_31_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_13_xor_79_nl = R_31_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_14_xor_79_nl = R_31_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_15_xor_79_nl = R_31_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign operator_8_false_1_mux1h_43_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_19_nl,
      loop_DES_rounds_4_xor_79_nl, loop_DES_rounds_5_xor_79_nl, loop_DES_rounds_6_xor_79_nl,
      loop_DES_rounds_7_xor_79_nl, loop_DES_rounds_8_xor_79_nl, loop_DES_rounds_9_xor_79_nl,
      loop_DES_rounds_10_xor_79_nl, loop_DES_rounds_11_xor_79_nl, loop_DES_rounds_12_xor_79_nl,
      loop_DES_rounds_13_xor_79_nl, loop_DES_rounds_14_xor_79_nl, loop_DES_rounds_15_xor_79_nl,
      loop_DES_rounds_8_xor_81, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_20_nl = (key_io_read_key_rsc_cse_63_1_sva[10]) ^ (reg_input_ftd[32])
      ^ (s_output_1_3_0_39_sva[2]);
  assign loop_DES_rounds_4_xor_75_nl = R_3_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_5_xor_75_nl = R_3_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_6_xor_75_nl = R_3_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_7_xor_75_nl = R_3_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_8_xor_75_nl = R_3_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_9_xor_75_nl = R_3_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_11_xor_75_nl = R_3_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_12_xor_75_nl = R_3_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_13_xor_75_nl = R_3_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_14_xor_75_nl = R_3_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_15_xor_75_nl = R_3_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_16_xor_75_nl = R_3_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign operator_8_false_1_mux1h_44_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_20_nl,
      loop_DES_rounds_4_xor_75_nl, loop_DES_rounds_5_xor_75_nl, loop_DES_rounds_6_xor_75_nl,
      loop_DES_rounds_7_xor_75_nl, loop_DES_rounds_8_xor_75_nl, loop_DES_rounds_9_xor_75_nl,
      loop_DES_rounds_4_xor_95, loop_DES_rounds_11_xor_75_nl, loop_DES_rounds_12_xor_75_nl,
      loop_DES_rounds_13_xor_75_nl, loop_DES_rounds_14_xor_75_nl, loop_DES_rounds_15_xor_75_nl,
      loop_DES_rounds_16_xor_75_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_21_nl = (reg_input_ftd[40]) ^ (s_output_1_19_16_50_sva[1])
      ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_4_xor_76_nl = R_2_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_5_xor_76_nl = R_1_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_6_xor_76_nl = R_10_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_7_xor_76_nl = R_20_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_8_xor_76_nl = R_11_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign loop_DES_rounds_9_xor_76_nl = R_31_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_10_xor_76_nl = R_2_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_11_xor_76_nl = R_19_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_12_xor_76_nl = R_1_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_13_xor_76_nl = R_19_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_14_xor_76_nl = R_10_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_15_xor_76_nl = R_19_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[34]);
  assign loop_DES_rounds_16_xor_76_nl = R_18_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign operator_8_false_1_mux1h_45_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_21_nl,
      loop_DES_rounds_4_xor_76_nl, loop_DES_rounds_5_xor_76_nl, loop_DES_rounds_6_xor_76_nl,
      loop_DES_rounds_7_xor_76_nl, loop_DES_rounds_8_xor_76_nl, loop_DES_rounds_9_xor_76_nl,
      loop_DES_rounds_10_xor_76_nl, loop_DES_rounds_11_xor_76_nl, loop_DES_rounds_12_xor_76_nl,
      loop_DES_rounds_13_xor_76_nl, loop_DES_rounds_14_xor_76_nl, loop_DES_rounds_15_xor_76_nl,
      loop_DES_rounds_16_xor_76_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_22_nl = (reg_input_ftd[48]) ^ (key_io_read_key_rsc_cse_63_1_sva[25])
      ^ (s_output_1_19_16_20_sva[0]);
  assign loop_DES_rounds_4_xor_77_nl = R_0_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_6_xor_77_nl = R_0_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_7_xor_77_nl = R_1_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_9_xor_77_nl = R_1_8_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_10_xor_77_nl = R_1_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[35]);
  assign loop_DES_rounds_11_xor_77_nl = R_0_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[51]);
  assign loop_DES_rounds_12_xor_77_nl = R_0_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign loop_DES_rounds_13_xor_77_nl = R_0_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_14_xor_77_nl = R_0_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_15_xor_77_nl = R_1_14_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_16_xor_77_nl = R_0_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign operator_8_false_1_mux1h_46_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_22_nl,
      loop_DES_rounds_4_xor_77_nl, loop_DES_rounds_5_xor_87, loop_DES_rounds_6_xor_77_nl,
      loop_DES_rounds_7_xor_77_nl, loop_DES_rounds_8_xor_87, loop_DES_rounds_9_xor_77_nl,
      loop_DES_rounds_10_xor_77_nl, loop_DES_rounds_11_xor_77_nl, loop_DES_rounds_12_xor_77_nl,
      loop_DES_rounds_13_xor_77_nl, loop_DES_rounds_14_xor_77_nl, loop_DES_rounds_15_xor_77_nl,
      loop_DES_rounds_16_xor_77_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign loop_DES_rounds_xor_23_nl = (reg_input_ftd[56]) ^ (s_output_1_3_0_54_sva[3])
      ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_4_xor_78_nl = R_0_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_5_xor_78_nl = R_0_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_6_xor_78_nl = R_0_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[17]);
  assign loop_DES_rounds_7_xor_78_nl = R_0_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_8_xor_78_nl = R_0_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_9_xor_78_nl = R_0_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_10_xor_78_nl = R_0_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[10]);
  assign loop_DES_rounds_11_xor_78_nl = R_0_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[26]);
  assign loop_DES_rounds_12_xor_78_nl = R_0_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_13_xor_78_nl = R_0_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_15_xor_78_nl = R_0_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_16_xor_78_nl = R_0_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[0]);
  assign operator_8_false_1_mux1h_47_nl = MUX1HOT_s_1_14_2(loop_DES_rounds_xor_23_nl,
      loop_DES_rounds_4_xor_78_nl, loop_DES_rounds_5_xor_78_nl, loop_DES_rounds_6_xor_78_nl,
      loop_DES_rounds_7_xor_78_nl, loop_DES_rounds_8_xor_78_nl, loop_DES_rounds_9_xor_78_nl,
      loop_DES_rounds_10_xor_78_nl, loop_DES_rounds_11_xor_78_nl, loop_DES_rounds_12_xor_78_nl,
      loop_DES_rounds_13_xor_78_nl, loop_DES_rounds_10_xor_85, loop_DES_rounds_15_xor_78_nl,
      loop_DES_rounds_16_xor_78_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])
      , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[15])});
  assign nl_U_ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_10_rg_I_1 = {operator_8_false_1_mux1h_7_nl
      , operator_8_false_1_mux1h_43_nl , operator_8_false_1_mux1h_44_nl , operator_8_false_1_mux1h_45_nl
      , operator_8_false_1_mux1h_46_nl , operator_8_false_1_mux1h_47_nl};
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd64)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd64)) key_rsci (
      .dat(key_rsc_dat),
      .idat(key_rsci_idat)
    );
  ccs_out_v1 #(.rscid(32'sd3),
  .width(32'sd64)) return_rsci (
      .idat(nl_return_rsci_idat[63:0]),
      .dat(return_rsc_dat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) input_rsc_triosy_obj (
      .ld(reg_key_rsc_triosy_obj_ld_cse),
      .lz(input_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) key_rsc_triosy_obj (
      .ld(reg_key_rsc_triosy_obj_ld_cse),
      .lz(key_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) return_rsc_triosy_obj (
      .ld(return_rsc_triosy_obj_ld),
      .lz(return_rsc_triosy_lz)
    );
  ROM_1i6_1o4_cfafff97e973ca9580e646fecdc2f814b3  U_ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_1_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_1_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_16)
    );
  ROM_1i6_1o4_d0e242163cbb0b2ce9c4399bc1cb50f5b3  U_ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_1_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_1_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_17)
    );
  ROM_1i6_1o4_752c7ca65a598ada4acee0cd63d199c3b3  U_ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_1_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_1_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_16)
    );
  ROM_1i6_1o4_ef717c7c87dc90ac6f7b34d533fe115fb3  U_ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_1_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_1_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_16)
    );
  ROM_1i6_1o4_3c5c29b75c561d2b741f22e5a3a569dbb3  U_ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_1_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_1_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_16)
    );
  ROM_1i6_1o4_ef4da7ff735c86ba85f23e51741d972cb3  U_ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_1_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_1_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_16)
    );
  ROM_1i6_1o4_ef4da7ff735c86ba85f23e51741d972cb3  U_ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_17)
    );
  ROM_1i6_1o4_752c7ca65a598ada4acee0cd63d199c3b3  U_ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_17)
    );
  ROM_1i6_1o4_3c5c29b75c561d2b741f22e5a3a569dbb3  U_ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_17)
    );
  ROM_1i6_1o4_51ba7157b272cd3b87451219caf38e7cb3  U_ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_17)
    );
  ROM_1i6_1o4_ef717c7c87dc90ac6f7b34d533fe115fb3  U_ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_17)
    );
  ROM_1i6_1o4_cfafff97e973ca9580e646fecdc2f814b3  U_ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_17)
    );
  ROM_1i6_1o4_cfafff97e973ca9580e646fecdc2f814b3  U_ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_10_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_10_rg_I_1[5:0]),
      .O_1(O_1_out)
    );
  ROM_1i6_1o4_d0e242163cbb0b2ce9c4399bc1cb50f5b3  U_ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_rg_I_1[5:0]),
      .O_1(O_1_out_1)
    );
  ROM_1i6_1o4_8f60b2fc4a3ee4cef30040071bc0219cb3  U_ROM_1i6_1o4_ce1b43b29576509b87f48de0e64c68b52f_1_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_ce1b43b29576509b87f48de0e64c68b52f_1_rg_I_1[5:0]),
      .O_1(O_1_out_2)
    );
  ROM_1i6_1o4_8f60b2fc4a3ee4cef30040071bc0219cb3  U_ROM_1i6_1o4_ce1b43b29576509b87f48de0e64c68b52f_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_ce1b43b29576509b87f48de0e64c68b52f_rg_I_1[5:0]),
      .O_1(O_1_out_3)
    );
  ROM_1i6_1o4_752c7ca65a598ada4acee0cd63d199c3b3  U_ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_10_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_10_rg_I_1[5:0]),
      .O_1(O_1_out_4)
    );
  ROM_1i6_1o4_ef717c7c87dc90ac6f7b34d533fe115fb3  U_ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_10_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_10_rg_I_1[5:0]),
      .O_1(O_1_out_5)
    );
  ROM_1i6_1o4_3c5c29b75c561d2b741f22e5a3a569dbb3  U_ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_10_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_10_rg_I_1[5:0]),
      .O_1(O_1_out_6)
    );
  ROM_1i6_1o4_51ba7157b272cd3b87451219caf38e7cb3  U_ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_1_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_1_rg_I_1[5:0]),
      .O_1(O_1_out_7)
    );
  ROM_1i6_1o4_ef4da7ff735c86ba85f23e51741d972cb3  U_ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_10_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_10_rg_I_1[5:0]),
      .O_1(O_1_out_8)
    );
  des_check_core_core_fsm des_check_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output)
    );
  assign loop_DES_rounds_16_xor_17_cse = R_7_1_sva ^ (O_1_out_5[1]);
  assign loop_DES_rounds_16_xor_32_cse = R_31_10_sva ^ (O_1_out_1[0]);
  assign loop_DES_rounds_16_xor_19_cse = R_30_4_sva ^ (O_1_out_1[3]);
  assign loop_DES_rounds_16_xor_14_cse = R_21_7_sva ^ (O_1_out_1[1]);
  assign loop_DES_rounds_16_xor_30_cse = R_3_4_sva ^ (O_1_out[1]);
  assign loop_DES_rounds_16_xor_21_cse = R_4_4_sva ^ (O_1_out_8[2]);
  assign loop_DES_rounds_16_xor_5_cse = R_12_4_sva ^ (O_1_out_7[0]);
  assign loop_DES_rounds_16_xor_12_cse = R_20_4_sva ^ (O_1_out_7[1]);
  assign loop_DES_rounds_16_xor_28_cse = R_28_4_sva ^ (O_1_out_5[0]);
  assign loop_DES_rounds_16_xor_23_cse = R_31_4_sva ^ (O_1_out[2]);
  assign loop_DES_rounds_16_xor_7_cse = R_11_4_sva ^ (O_1_out_1[2]);
  assign loop_DES_rounds_16_xor_10_cse = R_20_1_sva ^ (O_1_out_4[2]);
  assign loop_DES_rounds_16_xor_26_cse = R_27_4_sva ^ (O_1_out_7[3]);
  assign loop_DES_rounds_16_xor_25_cse = R_3_1_sva ^ (O_1_out_7[2]);
  assign loop_DES_rounds_16_xor_9_cse = R_11_1_sva ^ (O_1_out_8[0]);
  assign loop_DES_rounds_16_xor_8_cse = R_1_6_sva ^ (O_1_out[3]);
  assign loop_DES_rounds_16_xor_24_cse = R_27_10_sva ^ (O_1_out_8[3]);
  assign loop_DES_rounds_16_xor_27_cse = R_19_4_sva ^ (O_1_out_6[1]);
  assign loop_DES_rounds_16_xor_22_cse = R_25_6_sva ^ (O_1_out_6[0]);
  assign loop_DES_rounds_16_xor_4_cse = R_16_4_sva ^ (O_1_out_8[1]);
  assign loop_DES_rounds_16_xor_20_cse = R_24_4_sva ^ (O_1_out_4[0]);
  assign loop_DES_rounds_16_xor_31_cse = R_0_10_sva ^ (O_1_out_4[3]);
  assign loop_DES_rounds_16_xor_15_cse = R_7_4_sva ^ (O_1_out_6[3]);
  assign loop_DES_rounds_16_xor_2_cse = R_15_4_sva ^ (O_1_out_6[2]);
  assign loop_DES_rounds_16_xor_18_cse = R_23_4_sva ^ (O_1_out_5[3]);
  assign R_or_cse = (fsm_output[5]) | (fsm_output[7]);
  assign loop_DES_rounds_11_xor_13_cse = R_14_3_sva ^ (O_1_out_3[1]);
  assign loop_DES_rounds_6_xor_21_cse = R_0_1_sva ^ (O_1_out_8[2]);
  assign loop_DES_rounds_13_xor_13_cse = R_0_1_sva ^ (O_1_out_3[1]);
  assign R_or_1_cse = (fsm_output[0]) | (fsm_output[2]) | (fsm_output[4]) | (fsm_output[7])
      | (fsm_output[9]) | (fsm_output[11]) | (fsm_output[13]);
  assign R_or_133_cse = (fsm_output[11]) | (fsm_output[13]);
  assign loop_DES_rounds_5_xor_6_cse = R_18_3_sva ^ (O_1_out_5[2]);
  assign loop_DES_rounds_10_xor_25_cse = R_3_4_sva ^ (O_1_out_7[2]);
  assign R_or_2_cse = (fsm_output[0]) | (fsm_output[2]) | (fsm_output[4]) | (fsm_output[6])
      | (fsm_output[9]) | (fsm_output[11]) | (fsm_output[13]);
  assign loop_DES_rounds_10_xor_17_cse = R_7_4_sva ^ (O_1_out_5[1]);
  assign loop_DES_rounds_10_xor_14_cse = R_15_1_sva ^ (O_1_out_1[1]);
  assign loop_DES_rounds_5_xor_27_cse = R_2_3_sva ^ (O_1_out_6[1]);
  assign R_or_4_cse = (fsm_output[0]) | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[5])
      | (fsm_output[7]) | (fsm_output[9]) | (fsm_output[11]) | (fsm_output[13]);
  assign loop_DES_rounds_8_xor_4_cse = R_15_9_sva ^ (O_1_out_8[1]);
  assign loop_DES_rounds_10_xor_10_cse = R_20_4_sva ^ (O_1_out_4[2]);
  assign loop_DES_rounds_10_xor_9_cse = R_11_4_sva ^ (O_1_out_8[0]);
  assign R_or_127_cse = (fsm_output[12]) | (fsm_output[14]);
  assign loop_DES_rounds_11_xor_20_cse = R_24_11_sva ^ (O_1_out_4[0]);
  assign R_or_120_cse = (fsm_output[4]) | (fsm_output[6]) | (fsm_output[11]) | (fsm_output[13]);
  assign loop_DES_rounds_3_xor_31_cse = R_0_1_sva ^ (O_1_out_4[3]);
  assign loop_DES_rounds_10_xor_31_cse = R_0_4_sva ^ (O_1_out_4[3]);
  assign R_or_8_cse = (fsm_output[0]) | (fsm_output[2]) | (fsm_output[4]) | (fsm_output[6])
      | (fsm_output[8]) | (fsm_output[10]) | (fsm_output[12]) | (fsm_output[14]);
  assign R_or_122_cse = (fsm_output[4]) | (fsm_output[6]) | (fsm_output[8]);
  assign loop_DES_rounds_11_xor_9_cse = R_11_3_sva ^ (O_1_out_8[0]);
  assign loop_DES_rounds_5_xor_7_cse = R_11_11_sva ^ (O_1_out_1[2]);
  assign loop_DES_rounds_5_xor_1_cse = R_15_10_sva ^ (O_1_out_3[2]);
  assign loop_DES_rounds_3_xor_1_cse = R_15_1_sva ^ (O_1_out_3[2]);
  assign loop_DES_rounds_10_xor_1_cse = R_15_4_sva ^ (O_1_out_3[2]);
  assign loop_DES_rounds_11_xor_2_cse = R_16_3_sva ^ (O_1_out_6[2]);
  assign R_or_118_cse = (fsm_output[4]) | (fsm_output[6]) | (fsm_output[8]) | (fsm_output[10])
      | (fsm_output[12]) | (fsm_output[14]);
  assign loop_DES_rounds_6_xor_16_cse = R_23_4_sva ^ (O_1_out_3[3]);
  assign loop_DES_rounds_4_xor_16_cse = R_1_8_sva ^ (O_1_out_3[3]);
  assign loop_DES_rounds_10_xor_18_cse = R_24_4_sva ^ (O_1_out_5[3]);
  assign loop_DES_rounds_5_xor_18_cse = R_24_3_sva ^ (O_1_out_5[3]);
  assign loop_DES_rounds_15_xor_28_cse = R_26_4_sva ^ (O_1_out_5[0]);
  assign loop_DES_rounds_6_xor_24_cse = R_27_4_sva ^ (O_1_out_8[3]);
  assign loop_DES_rounds_10_xor_26_cse = R_28_4_sva ^ (O_1_out_7[3]);
  assign loop_DES_rounds_11_xor_32_cse = R_31_3_sva ^ (O_1_out_1[0]);
  assign loop_DES_rounds_5_xor_23_cse = R_31_11_sva ^ (O_1_out[2]);
  assign loop_DES_rounds_6_xor_32_cse = R_31_4_sva ^ (O_1_out_1[0]);
  assign loop_DES_rounds_10_xor_23_cse = R_4_4_sva ^ (O_1_out[2]);
  assign loop_DES_rounds_11_xor_17_cse = R_7_3_sva ^ (O_1_out_5[1]);
  assign loop_DES_rounds_5_xor_15_cse = R_7_11_sva ^ (O_1_out_6[3]);
  assign loop_DES_rounds_3_xor_15_cse = R_7_3_sva ^ (O_1_out_6[3]);
  assign loop_DES_rounds_5_xor_11_cse = R_10_10_sva ^ (O_1_out_4[1]);
  assign loop_DES_rounds_9_xor_5_cse = R_12_11_sva ^ (O_1_out_7[0]);
  assign loop_DES_rounds_5_xor_29_cse = R_0_11_sva ^ (O_1_out_3[0]);
  assign R_or_26_cse = (fsm_output[1]) | (fsm_output[2]) | (fsm_output[4]) | (fsm_output[6])
      | (fsm_output[8]) | (fsm_output[10]) | (fsm_output[12]);
  assign loop_DES_rounds_13_xor_4_cse = R_16_3_sva ^ (O_1_out_8[1]);
  assign loop_DES_rounds_11_xor_4_cse = R_15_11_sva ^ (O_1_out_8[1]);
  assign loop_DES_rounds_5_xor_25_cse = R_3_3_sva ^ (O_1_out_7[2]);
  assign loop_DES_rounds_4_xor_29_cse = R_0_4_sva ^ (O_1_out_3[0]);
  assign loop_DES_rounds_11_xor_11_cse = R_1_4_sva ^ (O_1_out_4[1]);
  assign loop_DES_rounds_10_xor_8_cse = R_19_4_sva ^ (O_1_out[3]);
  assign loop_DES_rounds_5_xor_12_cse = R_21_3_sva ^ (O_1_out_7[1]);
  assign R_or_32_cse = (fsm_output[2]) | (fsm_output[8]) | (fsm_output[10]) | (fsm_output[12])
      | (fsm_output[14]);
  assign loop_DES_rounds_11_xor_12_cse = R_21_7_sva ^ (O_1_out_7[1]);
  assign loop_DES_rounds_11_xor_14_cse = R_22_7_sva ^ (O_1_out_1[1]);
  assign R_or_105_cse = (fsm_output[6]) | (fsm_output[8]);
  assign loop_DES_rounds_15_xor_29_cse = R_0_9_sva ^ (O_1_out_3[0]);
  assign R_or_38_cse = (fsm_output[2]) | (fsm_output[3]) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[9]) | (fsm_output[11]) | (fsm_output[13]);
  assign loop_DES_rounds_10_xor_7_cse = R_12_4_sva ^ (O_1_out_1[2]);
  assign R_or_39_cse = (fsm_output[2]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[8])
      | (fsm_output[10]) | (fsm_output[12]) | (fsm_output[14]);
  assign loop_DES_rounds_10_xor_2_cse = R_16_4_sva ^ (O_1_out_6[2]);
  assign loop_DES_rounds_10_xor_20_cse = R_25_6_sva ^ (O_1_out_4[0]);
  assign loop_DES_rounds_10_xor_28_cse = R_29_4_sva ^ (O_1_out_5[0]);
  assign loop_DES_rounds_5_xor_30_cse = R_3_11_sva ^ (O_1_out[1]);
  assign loop_DES_rounds_10_xor_30_cse = R_30_4_sva ^ (O_1_out[1]);
  assign loop_DES_rounds_6_xor_6_cse = R_27_10_sva ^ (O_1_out_5[2]);
  assign loop_DES_rounds_4_xor_3_cse = R_1_14_sva ^ (O_1_out[0]);
  assign loop_DES_rounds_5_xor_21_cse = R_4_11_sva ^ (O_1_out_8[2]);
  assign loop_DES_rounds_10_xor_15_cse = R_8_4_sva ^ (O_1_out_6[3]);
  assign loop_DES_rounds_12_xor_13_cse = R_8_4_sva ^ (O_1_out_3[1]);
  assign loop_DES_rounds_10_xor_13_cse = R_9_4_sva ^ (O_1_out_3[1]);
  assign loop_DES_rounds_6_xor_19_cse = R_1_14_sva ^ (O_1_out_1[3]);
  assign loop_DES_rounds_10_xor_22_cse = R_26_4_sva ^ (O_1_out_6[0]);
  assign loop_DES_rounds_15_xor_21_cse = R_29_4_sva ^ (O_1_out_8[2]);
  assign loop_DES_rounds_13_xor_30_cse = R_26_5_sva ^ (O_1_out[1]);
  assign loop_DES_rounds_7_xor_22_cse = R_26_5_sva ^ (O_1_out_6[0]);
  assign loop_DES_rounds_13_xor_19_cse = R_29_5_sva ^ (O_1_out_1[3]);
  assign loop_DES_rounds_11_xor_19_cse = R_6_5_sva ^ (O_1_out_1[3]);
  assign loop_DES_rounds_7_xor_28_cse = R_29_5_sva ^ (O_1_out_5[0]);
  assign R_or_66_cse = (fsm_output[3]) | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[10])
      | (fsm_output[12]) | (fsm_output[14]);
  assign loop_DES_rounds_9_xor_81 = R_20_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[22]);
  assign loop_DES_rounds_5_xor_81 = R_15_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_7_xor_81 = R_7_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_8_xor_81 = R_31_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[24]);
  assign loop_DES_rounds_6_xor_81 = R_11_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[25]);
  assign loop_DES_rounds_9_xor_83 = R_27_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign loop_DES_rounds_8_xor_83 = R_24_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[28]);
  assign loop_DES_rounds_10_xor_81 = R_26_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[30]);
  assign loop_DES_rounds_8_xor_85 = R_11_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[32]);
  assign loop_DES_rounds_10_xor_83 = R_15_9_sva ^ (key_io_read_key_rsc_cse_63_1_sva[33]);
  assign loop_DES_rounds_4_xor_81 = R_25_6_sva ^ (key_io_read_key_rsc_cse_63_1_sva[36]);
  assign loop_DES_rounds_7_xor_83 = R_24_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[38]);
  assign loop_DES_rounds_4_xor_83 = R_4_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[40]);
  assign loop_DES_rounds_9_xor_85 = R_11_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[41]);
  assign loop_DES_rounds_4_xor_85 = R_7_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_8_xor_87 = R_1_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[42]);
  assign loop_DES_rounds_4_xor_87 = R_7_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_10_xor_85 = R_0_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[43]);
  assign loop_DES_rounds_2_xor_81 = R_23_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[44]);
  assign loop_DES_rounds_10_xor_87 = R_7_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_6_xor_83 = R_11_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[1]);
  assign loop_DES_rounds_4_xor_89 = R_29_5_sva ^ (key_io_read_key_rsc_cse_63_1_sva[2]);
  assign loop_DES_rounds_2_xor_83 = R_23_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[3]);
  assign loop_DES_rounds_2_xor_85 = R_7_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_9_xor_87 = R_7_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[48]);
  assign loop_DES_rounds_2_xor_87 = R_15_10_sva ^ (key_io_read_key_rsc_cse_63_1_sva[49]);
  assign loop_DES_rounds_8_xor_89 = R_12_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[50]);
  assign loop_DES_rounds_5_xor_83 = R_24_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[6]);
  assign loop_DES_rounds_10_xor_89 = R_24_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[52]);
  assign loop_DES_rounds_6_xor_85 = R_7_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[8]);
  assign loop_DES_rounds_7_xor_85 = R_28_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[53]);
  assign loop_DES_rounds_9_xor_89 = R_20_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[54]);
  assign loop_DES_rounds_2_xor_89 = R_28_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_6_xor_87 = R_20_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[11]);
  assign loop_DES_rounds_4_xor_91 = R_11_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign loop_DES_rounds_7_xor_87 = R_15_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[56]);
  assign loop_DES_rounds_4_xor_93 = R_21_7_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_5_xor_85 = R_23_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[12]);
  assign loop_DES_rounds_2_xor_91 = R_3_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_5_xor_87 = R_1_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[57]);
  assign loop_DES_rounds_9_xor_91 = R_3_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[58]);
  assign loop_DES_rounds_6_xor_89 = R_15_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[14]);
  assign loop_DES_rounds_5_xor_89 = R_7_4_sva ^ (key_io_read_key_rsc_cse_63_1_sva[59]);
  assign loop_DES_rounds_14_xor_81 = R_24_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[60]);
  assign loop_DES_rounds_4_xor_95 = R_3_3_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_2_xor_93 = R_0_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[16]);
  assign loop_DES_rounds_6_xor_91 = R_24_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_4_xor_97 = R_23_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[61]);
  assign loop_DES_rounds_2_xor_95 = R_7_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_6_xor_93 = R_12_11_sva ^ (key_io_read_key_rsc_cse_63_1_sva[18]);
  assign loop_DES_rounds_9_xor_93 = R_15_1_sva ^ (key_io_read_key_rsc_cse_63_1_sva[19]);
  always @(posedge clk) begin
    if ( rst ) begin
      key_io_read_key_rsc_cse_63_1_sva <= 63'b000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( fsm_output[0] ) begin
      key_io_read_key_rsc_cse_63_1_sva <= key_rsci_idat[63:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_0 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_0 <= loop_DES_rounds_16_xor_17_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_1 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_1 <= R_7_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_2 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_2 <= R_15_10_sva ^ (O_1_out_2[2]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_3 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_3 <= R_15_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_4 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_4 <= R_1_8_sva ^ (O_1_out_2[3]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_5 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_5 <= R_23_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_6 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_6 <= loop_DES_rounds_16_xor_32_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_7 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_7 <= R_31_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_8 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_8 <= loop_DES_rounds_16_xor_19_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_9 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_9 <= R_29_4_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_10 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_10 <= R_10_1_sva ^ (O_1_out[0]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_11 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_11 <= R_0_1_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_12 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_12 <= loop_DES_rounds_16_xor_14_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_13 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_13 <= R_21_3_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_14 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_14 <= loop_DES_rounds_16_xor_30_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_15 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_15 <= R_26_4_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_16 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_16 <= loop_DES_rounds_16_xor_21_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_17 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_17 <= R_26_5_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_18 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_18 <= loop_DES_rounds_16_xor_5_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_19 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_19 <= R_11_3_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_20 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_20 <= loop_DES_rounds_16_xor_12_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_21 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_21 <= R_2_3_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_22 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_22 <= loop_DES_rounds_16_xor_28_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_23 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_23 <= R_24_3_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_24 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_24 <= loop_DES_rounds_16_xor_23_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_25 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_25 <= R_4_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_26 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_26 <= loop_DES_rounds_16_xor_7_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_27 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_27 <= R_12_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_28 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_28 <= loop_DES_rounds_16_xor_10_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_29 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_29 <= R_20_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_30 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_30 <= loop_DES_rounds_16_xor_26_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_31 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_31 <= R_28_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_32 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_32 <= loop_DES_rounds_16_xor_25_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_33 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_33 <= R_3_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_34 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_34 <= loop_DES_rounds_16_xor_9_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_35 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_35 <= R_11_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_36 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_36 <= loop_DES_rounds_16_xor_8_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_37 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_37 <= R_19_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_38 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_38 <= loop_DES_rounds_16_xor_24_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_39 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_39 <= R_27_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_40 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_40 <= loop_DES_rounds_16_xor_27_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_41 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_41 <= R_18_3_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_42 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_42 <= R_1_7_sva ^ (O_1_out_4[1]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_43 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_43 <= R_0_9_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_44 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_44 <= R_31_3_sva ^ (O_1_out_5[2]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_45 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_45 <= R_1_4_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_46 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_46 <= loop_DES_rounds_16_xor_22_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_47 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_47 <= R_22_7_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_48 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_48 <= R_1_14_sva ^ (O_1_out_2[0]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_49 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_49 <= R_0_4_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_50 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_50 <= R_8_4_sva ^ (O_1_out_2[1]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_51 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_51 <= R_29_5_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_52 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_52 <= loop_DES_rounds_16_xor_4_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_53 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_53 <= R_14_3_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_54 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_54 <= loop_DES_rounds_16_xor_20_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_55 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_55 <= R_15_1_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_56 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_56 <= loop_DES_rounds_16_xor_31_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_57 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_57 <= R_0_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_58 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_58 <= loop_DES_rounds_16_xor_15_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_59 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_59 <= R_7_3_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_60 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_60 <= loop_DES_rounds_16_xor_2_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_61 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_61 <= R_15_9_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_62 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_62 <= loop_DES_rounds_16_xor_18_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_63 <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      return_rsci_idat_63 <= R_24_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_0_1_sva <= 1'b0;
    end
    else if ( (fsm_output[0]) | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[5])
        | (fsm_output[7]) | (fsm_output[10]) | (fsm_output[12]) | (fsm_output[14])
        ) begin
      R_0_1_sva <= MUX1HOT_s_1_7_2(loop_DES_rounds_1_xor_31_nl, loop_DES_rounds_2_xor_31_nl,
          loop_DES_rounds_16_xor_21_cse, loop_DES_rounds_6_xor_21_cse, loop_DES_rounds_11_xor_13_cse,
          loop_DES_rounds_13_xor_13_cse, loop_DES_rounds_15_xor_3_nl, {(fsm_output[0])
          , (fsm_output[2]) , (fsm_output[3]) , R_or_cse , (fsm_output[10]) , (fsm_output[12])
          , (fsm_output[14])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_3_1_sva <= 1'b0;
      R_10_1_sva <= 1'b0;
      R_1_8_sva <= 1'b0;
    end
    else if ( R_or_1_cse ) begin
      R_3_1_sva <= MUX1HOT_s_1_6_2(loop_DES_rounds_1_xor_25_nl, loop_DES_rounds_2_xor_25_nl,
          loop_DES_rounds_5_xor_6_cse, loop_DES_rounds_8_xor_5_nl, loop_DES_rounds_10_xor_25_cse,
          loop_DES_rounds_16_xor_25_cse, {(fsm_output[0]) , (fsm_output[2]) , (fsm_output[4])
          , (fsm_output[7]) , (fsm_output[9]) , R_or_133_cse});
      R_10_1_sva <= MUX1HOT_s_1_7_2(loop_DES_rounds_1_xor_11_nl, loop_DES_rounds_2_xor_19_nl,
          loop_DES_rounds_5_xor_27_cse, loop_DES_rounds_8_xor_11_nl, loop_DES_rounds_10_xor_14_cse,
          loop_DES_rounds_12_xor_6_nl, loop_DES_rounds_14_xor_3_nl, {(fsm_output[0])
          , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])
          , (fsm_output[11]) , (fsm_output[13])});
      R_1_8_sva <= MUX1HOT_s_1_6_2(loop_DES_rounds_1_xor_22_nl, loop_DES_rounds_2_xor_16_nl,
          loop_DES_rounds_5_xor_11_cse, loop_DES_rounds_8_xor_29_nl, loop_DES_rounds_6_xor_16_cse,
          loop_DES_rounds_4_xor_16_cse, {(fsm_output[0]) , (fsm_output[2]) , (fsm_output[4])
          , (fsm_output[7]) , (fsm_output[9]) , R_or_133_cse});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_7_1_sva <= 1'b0;
      R_0_10_sva <= 1'b0;
      R_15_10_sva <= 1'b0;
    end
    else if ( R_or_2_cse ) begin
      R_7_1_sva <= MUX1HOT_s_1_6_2(loop_DES_rounds_1_xor_17_nl, loop_DES_rounds_2_xor_17_nl,
          loop_DES_rounds_5_xor_3_nl, loop_DES_rounds_7_xor_6_nl, loop_DES_rounds_10_xor_17_cse,
          loop_DES_rounds_16_xor_17_cse, {(fsm_output[0]) , (fsm_output[2]) , (fsm_output[4])
          , (fsm_output[6]) , (fsm_output[9]) , R_or_133_cse});
      R_0_10_sva <= MUX1HOT_s_1_4_2(loop_DES_rounds_1_xor_29_nl, loop_DES_rounds_3_xor_31_cse,
          loop_DES_rounds_16_xor_31_cse, loop_DES_rounds_10_xor_31_cse, {(fsm_output[0])
          , (fsm_output[2]) , R_or_120_cse , (fsm_output[9])});
      R_15_10_sva <= MUX1HOT_s_1_4_2(loop_DES_rounds_1_xor_2_nl, loop_DES_rounds_3_xor_1_cse,
          loop_DES_rounds_5_xor_1_cse, loop_DES_rounds_10_xor_1_cse, {(fsm_output[0])
          , (fsm_output[2]) , R_or_120_cse , (fsm_output[9])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_20_1_sva <= 1'b0;
      R_23_4_sva <= 1'b0;
      R_27_4_sva <= 1'b0;
      R_31_4_sva <= 1'b0;
    end
    else if ( R_or_4_cse ) begin
      R_20_1_sva <= MUX1HOT_s_1_7_2(loop_DES_rounds_1_xor_10_nl, loop_DES_rounds_2_xor_10_nl,
          loop_DES_rounds_16_xor_5_cse, loop_DES_rounds_6_xor_27_nl, loop_DES_rounds_8_xor_4_cse,
          loop_DES_rounds_10_xor_10_cse, loop_DES_rounds_16_xor_10_cse, {(fsm_output[0])
          , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[7])
          , (fsm_output[9]) , R_or_133_cse});
      R_23_4_sva <= MUX1HOT_s_1_6_2(loop_DES_rounds_1_xor_4_nl, loop_DES_rounds_2_xor_18_nl,
          loop_DES_rounds_4_xor_16_cse, loop_DES_rounds_6_xor_16_cse, loop_DES_rounds_10_xor_18_cse,
          loop_DES_rounds_16_xor_18_cse, {(fsm_output[0]) , (fsm_output[2]) , (fsm_output[3])
          , R_or_cse , (fsm_output[9]) , R_or_133_cse});
      R_27_4_sva <= MUX1HOT_s_1_6_2(loop_DES_rounds_1_xor_6_nl, loop_DES_rounds_2_xor_26_nl,
          loop_DES_rounds_16_xor_24_cse, loop_DES_rounds_6_xor_24_cse, loop_DES_rounds_10_xor_26_cse,
          loop_DES_rounds_16_xor_26_cse, {(fsm_output[0]) , (fsm_output[2]) , (fsm_output[3])
          , R_or_cse , (fsm_output[9]) , R_or_133_cse});
      R_31_4_sva <= MUX1HOT_s_1_6_2(loop_DES_rounds_1_xor_24_nl, loop_DES_rounds_2_xor_23_nl,
          loop_DES_rounds_16_xor_32_cse, loop_DES_rounds_6_xor_32_cse, loop_DES_rounds_10_xor_23_cse,
          loop_DES_rounds_16_xor_23_cse, {(fsm_output[0]) , (fsm_output[2]) , (fsm_output[3])
          , R_or_cse , (fsm_output[9]) , R_or_133_cse});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_11_1_sva <= 1'b0;
    end
    else if ( (fsm_output[0]) | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6])
        | (fsm_output[9]) | (fsm_output[11]) | (fsm_output[13]) ) begin
      R_11_1_sva <= MUX1HOT_s_1_6_2(loop_DES_rounds_1_xor_9_nl, loop_DES_rounds_2_xor_9_nl,
          loop_DES_rounds_4_xor_14_nl, loop_DES_rounds_7_xor_27_nl, loop_DES_rounds_10_xor_9_cse,
          loop_DES_rounds_16_xor_9_cse, {(fsm_output[0]) , (fsm_output[2]) , (fsm_output[3])
          , (fsm_output[6]) , (fsm_output[9]) , R_or_133_cse});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_15_1_sva <= 1'b0;
    end
    else if ( (fsm_output[0]) | (fsm_output[2]) | (fsm_output[5]) | (fsm_output[7])
        | (fsm_output[10]) | (fsm_output[12]) | (fsm_output[14]) ) begin
      R_15_1_sva <= MUX1HOT_s_1_6_2(loop_DES_rounds_1_xor_1_nl, loop_DES_rounds_2_xor_1_nl,
          loop_DES_rounds_6_xor_14_nl, loop_DES_rounds_10_xor_14_cse, loop_DES_rounds_11_xor_20_cse,
          loop_DES_rounds_13_xor_20_nl, {(fsm_output[0]) , (fsm_output[2]) , (fsm_output[5])
          , (fsm_output[7]) , (fsm_output[10]) , R_or_127_cse});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      s_output_1_19_16_35_sva <= 4'b0000;
    end
    else if ( fsm_output[0] ) begin
      s_output_1_19_16_35_sva <= ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_16;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsc_triosy_obj_ld <= 1'b0;
      reg_key_rsc_triosy_obj_ld_cse <= 1'b0;
      s_output_1_19_16_20_sva <= 4'b0000;
      s_output_1_19_16_5_sva <= 4'b0000;
      s_output_1_3_0_54_sva <= 4'b0000;
      s_output_1_3_0_24_sva <= 4'b0000;
      s_output_1_19_16_50_sva <= 4'b0000;
      s_output_1_3_0_39_sva <= 4'b0000;
      s_output_1_3_0_9_sva <= 4'b0000;
    end
    else begin
      return_rsc_triosy_obj_ld <= fsm_output[15];
      reg_key_rsc_triosy_obj_ld_cse <= fsm_output[0];
      s_output_1_19_16_20_sva <= MUX_v_4_2_2(O_1_out_1, O_1_out_2, fsm_output[1]);
      s_output_1_19_16_5_sva <= ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_17;
      s_output_1_3_0_54_sva <= ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_16;
      s_output_1_3_0_24_sva <= ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_16;
      s_output_1_19_16_50_sva <= ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_16;
      s_output_1_3_0_39_sva <= O_1_out_7;
      s_output_1_3_0_9_sva <= ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_16;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_11_11_sva <= 1'b0;
      R_19_11_sva <= 1'b0;
      R_20_11_sva <= 1'b0;
      R_23_11_sva <= 1'b0;
      R_24_3_sva <= 1'b0;
      R_27_11_sva <= 1'b0;
      R_28_11_sva <= 1'b0;
      R_31_11_sva <= 1'b0;
      R_7_11_sva <= 1'b0;
      R_7_3_sva <= 1'b0;
    end
    else if ( R_or_8_cse ) begin
      R_11_11_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_1_xor_5_nl, loop_DES_rounds_3_xor_7_nl,
          loop_DES_rounds_5_xor_7_cse, loop_DES_rounds_11_xor_9_cse, loop_DES_rounds_13_xor_9_nl,
          {(fsm_output[0]) , (fsm_output[2]) , R_or_122_cse , (fsm_output[10]) ,
          R_or_127_cse});
      R_19_11_sva <= MUX1HOT_s_1_3_2(loop_DES_rounds_1_xor_27_nl, loop_DES_rounds_3_xor_8_nl,
          loop_DES_rounds_5_xor_8_nl, {(fsm_output[0]) , (fsm_output[2]) , R_or_118_cse});
      R_20_11_sva <= MUX1HOT_s_1_3_2(loop_DES_rounds_1_xor_12_nl, loop_DES_rounds_16_xor_10_cse,
          loop_DES_rounds_5_xor_10_nl, {(fsm_output[0]) , (fsm_output[2]) , R_or_118_cse});
      R_23_11_sva <= MUX1HOT_s_1_3_2(loop_DES_rounds_1_xor_18_nl, loop_DES_rounds_3_xor_16_nl,
          loop_DES_rounds_5_xor_16_nl, {(fsm_output[0]) , (fsm_output[2]) , R_or_118_cse});
      R_24_3_sva <= MUX1HOT_s_1_6_2(loop_DES_rounds_1_xor_20_nl, loop_DES_rounds_3_xor_18_nl,
          loop_DES_rounds_5_xor_18_cse, loop_DES_rounds_11_xor_5_nl, loop_DES_rounds_13_xor_6_nl,
          loop_DES_rounds_15_xor_28_cse, {(fsm_output[0]) , (fsm_output[2]) , R_or_122_cse
          , (fsm_output[10]) , (fsm_output[12]) , (fsm_output[14])});
      R_27_11_sva <= MUX1HOT_s_1_3_2(loop_DES_rounds_1_xor_26_nl, loop_DES_rounds_3_xor_24_nl,
          loop_DES_rounds_5_xor_24_nl, {(fsm_output[0]) , (fsm_output[2]) , R_or_118_cse});
      R_28_11_sva <= MUX1HOT_s_1_3_2(loop_DES_rounds_1_xor_28_nl, loop_DES_rounds_3_xor_26_nl,
          loop_DES_rounds_5_xor_26_nl, {(fsm_output[0]) , (fsm_output[2]) , R_or_118_cse});
      R_31_11_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_1_xor_21_nl, loop_DES_rounds_3_xor_23_nl,
          loop_DES_rounds_5_xor_23_cse, loop_DES_rounds_11_xor_32_cse, loop_DES_rounds_13_xor_32_nl,
          {(fsm_output[0]) , (fsm_output[2]) , R_or_122_cse , (fsm_output[10]) ,
          R_or_127_cse});
      R_7_11_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_1_xor_13_nl, loop_DES_rounds_3_xor_15_cse,
          loop_DES_rounds_5_xor_15_cse, loop_DES_rounds_11_xor_17_cse, loop_DES_rounds_13_xor_17_nl,
          {(fsm_output[0]) , (fsm_output[2]) , R_or_122_cse , (fsm_output[10]) ,
          R_or_127_cse});
      R_7_3_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_1_xor_15_nl, loop_DES_rounds_16_xor_17_cse,
          loop_DES_rounds_11_xor_17_cse, loop_DES_rounds_5_xor_15_cse, loop_DES_rounds_3_xor_15_cse,
          {(fsm_output[0]) , (fsm_output[2]) , R_or_122_cse , (fsm_output[10]) ,
          R_or_127_cse});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_15_9_sva <= 1'b0;
    end
    else if ( (fsm_output[3]) | (fsm_output[14]) | (fsm_output[0]) | (fsm_output[5])
        | (fsm_output[8]) | (fsm_output[10]) | (fsm_output[12]) ) begin
      R_15_9_sva <= MUX1HOT_s_1_6_2(loop_DES_rounds_1_xor_16_nl, loop_DES_rounds_16_xor_4_cse,
          loop_DES_rounds_8_xor_4_cse, loop_DES_rounds_5_xor_1_cse, loop_DES_rounds_11_xor_2_cse,
          loop_DES_rounds_13_xor_2_nl, {(fsm_output[0]) , (fsm_output[3]) , (fsm_output[5])
          , (fsm_output[8]) , (fsm_output[10]) , R_or_127_cse});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_0_11_sva <= 1'b0;
    end
    else if ( (fsm_output[1]) | (fsm_output[2]) | (fsm_output[4]) | (fsm_output[6])
        | (fsm_output[8]) | (fsm_output[10]) | (fsm_output[12]) | (fsm_output[14])
        ) begin
      R_0_11_sva <= MUX1HOT_s_1_7_2(loop_DES_rounds_1_xor_3_nl, loop_DES_rounds_3_xor_29_nl,
          loop_DES_rounds_5_xor_29_cse, loop_DES_rounds_7_xor_11_nl, loop_DES_rounds_9_xor_5_cse,
          loop_DES_rounds_11_xor_31_nl, loop_DES_rounds_13_xor_31_nl, {(fsm_output[1])
          , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])
          , (fsm_output[10]) , R_or_127_cse});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_11_3_sva <= 1'b0;
    end
    else if ( (fsm_output[1]) | (fsm_output[2]) | (fsm_output[4]) | (fsm_output[6])
        | (fsm_output[8]) | (fsm_output[14]) ) begin
      R_11_3_sva <= MUX1HOT_s_1_4_2(loop_DES_rounds_1_xor_7_nl, loop_DES_rounds_16_xor_9_cse,
          loop_DES_rounds_11_xor_9_cse, loop_DES_rounds_15_xor_5_nl, {(fsm_output[1])
          , (fsm_output[2]) , R_or_122_cse , (fsm_output[14])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_16_3_sva <= 1'b0;
      R_3_3_sva <= 1'b0;
    end
    else if ( R_or_26_cse ) begin
      R_16_3_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_1_xor_8_nl, loop_DES_rounds_3_xor_2_nl,
          loop_DES_rounds_11_xor_2_cse, loop_DES_rounds_11_xor_4_cse, loop_DES_rounds_13_xor_4_cse,
          {(fsm_output[1]) , (fsm_output[2]) , R_or_122_cse , (fsm_output[10]) ,
          (fsm_output[12])});
      R_3_3_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_1_xor_30_nl, loop_DES_rounds_16_xor_25_cse,
          loop_DES_rounds_5_xor_25_cse, loop_DES_rounds_5_xor_6_cse, loop_DES_rounds_13_xor_5_nl,
          {(fsm_output[1]) , (fsm_output[2]) , R_or_122_cse , (fsm_output[10]) ,
          (fsm_output[12])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_31_3_sva <= 1'b0;
    end
    else if ( (fsm_output[1]) | (fsm_output[2]) | (fsm_output[4]) | (fsm_output[6])
        | (fsm_output[8]) | (fsm_output[10]) | (fsm_output[13]) ) begin
      R_31_3_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_1_xor_23_nl, loop_DES_rounds_3_xor_32_nl,
          loop_DES_rounds_11_xor_32_cse, loop_DES_rounds_11_xor_3_nl, loop_DES_rounds_14_xor_6_nl,
          {(fsm_output[1]) , (fsm_output[2]) , R_or_122_cse , (fsm_output[10]) ,
          (fsm_output[13])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_1_4_sva <= 1'b0;
    end
    else if ( (fsm_output[1]) | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[5])
        | (fsm_output[8]) | (fsm_output[10]) | (fsm_output[12]) | (fsm_output[14])
        ) begin
      R_1_4_sva <= MUX1HOT_s_1_7_2(loop_DES_rounds_1_xor_19_nl, loop_DES_rounds_2_xor_6_nl,
          loop_DES_rounds_4_xor_29_cse, loop_DES_rounds_6_xor_3_nl, loop_DES_rounds_9_xor_11_nl,
          loop_DES_rounds_11_xor_11_cse, loop_DES_rounds_15_xor_6_nl, {(fsm_output[1])
          , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[8])
          , R_or_125_nl , (fsm_output[14])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_1_6_sva <= 1'b0;
    end
    else if ( (fsm_output[1]) | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[5])
        | (fsm_output[7]) | (fsm_output[9]) | (fsm_output[11]) | (fsm_output[13])
        ) begin
      R_1_6_sva <= MUX1HOT_s_1_7_2(loop_DES_rounds_1_xor_14_nl, loop_DES_rounds_2_xor_8_nl,
          loop_DES_rounds_4_xor_11_nl, loop_DES_rounds_6_xor_29_nl, loop_DES_rounds_8_xor_3_nl,
          loop_DES_rounds_10_xor_8_cse, loop_DES_rounds_16_xor_8_cse, {(fsm_output[1])
          , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[7])
          , (fsm_output[9]) , R_or_133_cse});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_10_10_sva <= 1'b0;
    end
    else if ( (fsm_output[12]) | (fsm_output[9]) | (fsm_output[6]) | (fsm_output[1])
        | (fsm_output[2]) | (fsm_output[4]) ) begin
      R_10_10_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_1_xor_32_nl, loop_DES_rounds_3_xor_11_nl,
          loop_DES_rounds_5_xor_12_cse, loop_DES_rounds_7_xor_3_nl, loop_DES_rounds_13_xor_27_nl,
          {(fsm_output[1]) , R_or_102_nl , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[12])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_2_3_sva <= 1'b0;
      R_0_9_sva <= 1'b0;
    end
    else if ( R_or_32_cse ) begin
      R_2_3_sva <= MUX1HOT_s_1_4_2(loop_DES_rounds_3_xor_27_nl, loop_DES_rounds_9_xor_27_nl,
          loop_DES_rounds_11_xor_12_cse, loop_DES_rounds_13_xor_12_nl, {(fsm_output[2])
          , (fsm_output[8]) , (fsm_output[10]) , R_or_127_cse});
      R_0_9_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_2_xor_11_nl, loop_DES_rounds_16_xor_31_cse,
          loop_DES_rounds_11_xor_29_nl, loop_DES_rounds_15_xor_29_cse, loop_DES_rounds_11_xor_11_cse,
          {(fsm_output[2]) , (fsm_output[8]) , (fsm_output[10]) , (fsm_output[12])
          , (fsm_output[14])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_21_3_sva <= 1'b0;
    end
    else if ( (fsm_output[5]) | (fsm_output[2]) | (fsm_output[14]) | (fsm_output[7])
        | (fsm_output[10]) | (fsm_output[12]) ) begin
      R_21_3_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_3_xor_12_nl, loop_DES_rounds_6_xor_12_nl,
          loop_DES_rounds_5_xor_12_cse, loop_DES_rounds_11_xor_14_cse, loop_DES_rounds_13_xor_14_nl,
          {(fsm_output[2]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[10])
          , R_or_127_cse});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_18_3_sva <= 1'b0;
    end
    else if ( (fsm_output[8]) | (fsm_output[2]) | (fsm_output[14]) ) begin
      R_18_3_sva <= MUX1HOT_s_1_3_2(loop_DES_rounds_3_xor_6_nl, loop_DES_rounds_9_xor_6_nl,
          loop_DES_rounds_15_xor_27_nl, {(fsm_output[2]) , (fsm_output[8]) , (fsm_output[14])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_14_3_sva <= 1'b0;
    end
    else if ( (fsm_output[2]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[8])
        | (fsm_output[14]) ) begin
      R_14_3_sva <= MUX1HOT_s_1_4_2(loop_DES_rounds_3_xor_3_nl, loop_DES_rounds_5_xor_13_nl,
          loop_DES_rounds_11_xor_13_cse, loop_DES_rounds_13_xor_4_cse, {(fsm_output[2])
          , (fsm_output[4]) , R_or_105_cse , (fsm_output[14])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_0_4_sva <= 1'b0;
    end
    else if ( (fsm_output[2]) | (fsm_output[3]) | (fsm_output[5]) | (fsm_output[7])
        | (fsm_output[9]) | (fsm_output[11]) | (fsm_output[14]) ) begin
      R_0_4_sva <= MUX1HOT_s_1_6_2(loop_DES_rounds_2_xor_29_nl, loop_DES_rounds_3_xor_31_cse,
          loop_DES_rounds_10_xor_31_cse, loop_DES_rounds_10_xor_29_nl, loop_DES_rounds_4_xor_29_cse,
          loop_DES_rounds_15_xor_29_cse, {(fsm_output[2]) , (fsm_output[3]) , R_or_cse
          , (fsm_output[9]) , (fsm_output[11]) , (fsm_output[14])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_11_4_sva <= 1'b0;
      R_12_4_sva <= 1'b0;
      R_15_4_sva <= 1'b0;
      R_16_4_sva <= 1'b0;
      R_19_4_sva <= 1'b0;
      R_20_4_sva <= 1'b0;
      R_24_4_sva <= 1'b0;
      R_27_10_sva <= 1'b0;
      R_28_4_sva <= 1'b0;
      R_3_4_sva <= 1'b0;
      R_31_10_sva <= 1'b0;
      R_4_4_sva <= 1'b0;
      R_7_4_sva <= 1'b0;
      R_8_4_sva <= 1'b0;
      R_1_14_sva <= 1'b0;
    end
    else if ( R_or_38_cse ) begin
      R_11_4_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_2_xor_7_nl, loop_DES_rounds_16_xor_9_cse,
          loop_DES_rounds_10_xor_9_cse, loop_DES_rounds_10_xor_7_cse, loop_DES_rounds_16_xor_7_cse,
          {(fsm_output[2]) , (fsm_output[3]) , R_or_cse , (fsm_output[9]) , R_or_133_cse});
      R_12_4_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_2_xor_5_nl, loop_DES_rounds_16_xor_7_cse,
          loop_DES_rounds_10_xor_7_cse, loop_DES_rounds_10_xor_5_nl, loop_DES_rounds_16_xor_5_cse,
          {(fsm_output[2]) , (fsm_output[3]) , R_or_cse , (fsm_output[9]) , R_or_133_cse});
      R_15_4_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_2_xor_2_nl, loop_DES_rounds_3_xor_1_cse,
          loop_DES_rounds_10_xor_1_cse, loop_DES_rounds_10_xor_2_cse, loop_DES_rounds_16_xor_2_cse,
          {(fsm_output[2]) , (fsm_output[3]) , R_or_cse , (fsm_output[9]) , R_or_133_cse});
      R_16_4_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_2_xor_4_nl, loop_DES_rounds_16_xor_2_cse,
          loop_DES_rounds_10_xor_2_cse, loop_DES_rounds_10_xor_4_nl, loop_DES_rounds_16_xor_4_cse,
          {(fsm_output[2]) , (fsm_output[3]) , R_or_cse , (fsm_output[9]) , R_or_133_cse});
      R_19_4_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_2_xor_27_nl, loop_DES_rounds_16_xor_8_cse,
          loop_DES_rounds_10_xor_8_cse, loop_DES_rounds_10_xor_27_nl, loop_DES_rounds_16_xor_27_cse,
          {(fsm_output[2]) , (fsm_output[3]) , R_or_cse , (fsm_output[9]) , R_or_133_cse});
      R_20_4_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_2_xor_12_nl, loop_DES_rounds_16_xor_10_cse,
          loop_DES_rounds_10_xor_10_cse, loop_DES_rounds_5_xor_12_cse, loop_DES_rounds_16_xor_12_cse,
          {(fsm_output[2]) , (fsm_output[3]) , R_or_cse , (fsm_output[9]) , R_or_133_cse});
      R_24_4_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_2_xor_20_nl, loop_DES_rounds_16_xor_18_cse,
          loop_DES_rounds_10_xor_18_cse, loop_DES_rounds_10_xor_20_cse, loop_DES_rounds_16_xor_20_cse,
          {(fsm_output[2]) , (fsm_output[3]) , R_or_cse , (fsm_output[9]) , R_or_133_cse});
      R_27_10_sva <= MUX1HOT_s_1_6_2(loop_DES_rounds_2_xor_24_nl, loop_DES_rounds_4_xor_6_nl,
          loop_DES_rounds_6_xor_5_nl, loop_DES_rounds_8_xor_6_nl, loop_DES_rounds_6_xor_24_cse,
          loop_DES_rounds_16_xor_24_cse, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[5])
          , (fsm_output[7]) , (fsm_output[9]) , R_or_133_cse});
      R_28_4_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_2_xor_28_nl, loop_DES_rounds_16_xor_26_cse,
          loop_DES_rounds_10_xor_26_cse, loop_DES_rounds_10_xor_28_cse, loop_DES_rounds_16_xor_28_cse,
          {(fsm_output[2]) , (fsm_output[3]) , R_or_cse , (fsm_output[9]) , R_or_133_cse});
      R_3_4_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_2_xor_30_nl, loop_DES_rounds_16_xor_25_cse,
          loop_DES_rounds_10_xor_25_cse, loop_DES_rounds_10_xor_30_cse, loop_DES_rounds_16_xor_30_cse,
          {(fsm_output[2]) , (fsm_output[3]) , R_or_cse , (fsm_output[9]) , R_or_133_cse});
      R_31_10_sva <= MUX1HOT_s_1_6_2(loop_DES_rounds_2_xor_32_nl, loop_DES_rounds_4_xor_3_cse,
          loop_DES_rounds_6_xor_6_cse, loop_DES_rounds_8_xor_27_nl, loop_DES_rounds_6_xor_32_cse,
          loop_DES_rounds_16_xor_32_cse, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[5])
          , (fsm_output[7]) , (fsm_output[9]) , R_or_133_cse});
      R_4_4_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_2_xor_21_nl, loop_DES_rounds_16_xor_23_cse,
          loop_DES_rounds_10_xor_23_cse, loop_DES_rounds_6_xor_21_cse, loop_DES_rounds_16_xor_21_cse,
          {(fsm_output[2]) , (fsm_output[3]) , R_or_cse , (fsm_output[9]) , R_or_133_cse});
      R_7_4_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_2_xor_15_nl, loop_DES_rounds_16_xor_17_cse,
          loop_DES_rounds_10_xor_17_cse, loop_DES_rounds_10_xor_15_cse, loop_DES_rounds_16_xor_15_cse,
          {(fsm_output[2]) , (fsm_output[3]) , R_or_cse , (fsm_output[9]) , R_or_133_cse});
      R_8_4_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_2_xor_13_nl, loop_DES_rounds_16_xor_15_cse,
          loop_DES_rounds_10_xor_15_cse, loop_DES_rounds_10_xor_13_cse, loop_DES_rounds_12_xor_13_cse,
          {(fsm_output[2]) , (fsm_output[3]) , R_or_cse , (fsm_output[9]) , R_or_133_cse});
      R_1_14_sva <= MUX1HOT_s_1_6_2(loop_DES_rounds_2_xor_3_nl, loop_DES_rounds_4_xor_19_nl,
          loop_DES_rounds_6_xor_19_cse, loop_DES_rounds_10_xor_3_nl, loop_DES_rounds_5_xor_11_cse,
          loop_DES_rounds_4_xor_29_cse, {(fsm_output[2]) , (fsm_output[3]) , R_or_cse
          , (fsm_output[9]) , (fsm_output[11]) , (fsm_output[13])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_12_11_sva <= 1'b0;
      R_15_11_sva <= 1'b0;
      R_24_11_sva <= 1'b0;
      R_3_11_sva <= 1'b0;
      R_4_11_sva <= 1'b0;
      R_26_5_sva <= 1'b0;
      R_29_5_sva <= 1'b0;
    end
    else if ( R_or_39_cse ) begin
      R_12_11_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_3_xor_5_nl, loop_DES_rounds_9_xor_5_cse,
          loop_DES_rounds_9_xor_3_nl, loop_DES_rounds_5_xor_7_cse, loop_DES_rounds_13_xor_7_nl,
          {(fsm_output[2]) , R_or_99_nl , (fsm_output[8]) , (fsm_output[10]) , R_or_127_cse});
      R_15_11_sva <= MUX1HOT_s_1_4_2(loop_DES_rounds_3_xor_4_nl, loop_DES_rounds_11_xor_4_cse,
          loop_DES_rounds_11_xor_1_nl, loop_DES_rounds_13_xor_1_nl, {(fsm_output[2])
          , R_or_122_cse , (fsm_output[10]) , R_or_127_cse});
      R_24_11_sva <= MUX1HOT_s_1_4_2(loop_DES_rounds_3_xor_20_nl, loop_DES_rounds_11_xor_20_cse,
          loop_DES_rounds_5_xor_18_cse, loop_DES_rounds_13_xor_18_nl, {(fsm_output[2])
          , R_or_122_cse , (fsm_output[10]) , R_or_127_cse});
      R_3_11_sva <= MUX1HOT_s_1_4_2(loop_DES_rounds_3_xor_30_nl, loop_DES_rounds_5_xor_30_cse,
          loop_DES_rounds_5_xor_25_cse, loop_DES_rounds_13_xor_25_nl, {(fsm_output[2])
          , R_or_122_cse , (fsm_output[10]) , R_or_127_cse});
      R_4_11_sva <= MUX1HOT_s_1_4_2(loop_DES_rounds_3_xor_21_nl, loop_DES_rounds_5_xor_21_cse,
          loop_DES_rounds_5_xor_23_cse, loop_DES_rounds_13_xor_23_nl, {(fsm_output[2])
          , R_or_122_cse , (fsm_output[10]) , R_or_127_cse});
      R_26_5_sva <= MUX1HOT_s_1_6_2(loop_DES_rounds_3_xor_28_nl, loop_DES_rounds_16_xor_22_cse,
          loop_DES_rounds_7_xor_22_cse, loop_DES_rounds_5_xor_30_cse, loop_DES_rounds_13_xor_30_cse,
          loop_DES_rounds_15_xor_21_cse, {(fsm_output[2]) , (fsm_output[4]) , R_or_105_cse
          , (fsm_output[10]) , (fsm_output[12]) , (fsm_output[14])});
      R_29_5_sva <= MUX1HOT_s_1_6_2(loop_DES_rounds_3_xor_19_nl, loop_DES_rounds_5_xor_28_nl,
          loop_DES_rounds_7_xor_28_cse, loop_DES_rounds_11_xor_19_cse, loop_DES_rounds_13_xor_19_cse,
          loop_DES_rounds_13_xor_13_cse, {(fsm_output[2]) , (fsm_output[4]) , R_or_105_cse
          , (fsm_output[10]) , (fsm_output[12]) , (fsm_output[14])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_1_7_sva <= 1'b0;
    end
    else if ( (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9])
        | (fsm_output[11]) | (fsm_output[13]) ) begin
      R_1_7_sva <= MUX1HOT_s_1_6_2(loop_DES_rounds_2_xor_14_nl, loop_DES_rounds_16_xor_27_cse,
          loop_DES_rounds_5_xor_29_cse, loop_DES_rounds_6_xor_6_cse, loop_DES_rounds_4_xor_3_cse,
          loop_DES_rounds_14_xor_11_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[6])
          , (fsm_output[9]) , (fsm_output[11]) , (fsm_output[13])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_1_9_sva <= 1'b0;
    end
    else if ( (fsm_output[2]) | (fsm_output[3]) | (fsm_output[5]) | (fsm_output[8])
        | (fsm_output[10]) | (fsm_output[12]) ) begin
      R_1_9_sva <= MUX1HOT_s_1_6_2(loop_DES_rounds_2_xor_22_nl, loop_DES_rounds_16_xor_12_cse,
          loop_DES_rounds_6_xor_11_nl, loop_DES_rounds_9_xor_29_nl, loop_DES_rounds_5_xor_27_cse,
          loop_DES_rounds_13_xor_3_nl, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[5])
          , (fsm_output[8]) , (fsm_output[10]) , (fsm_output[12])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_21_7_sva <= 1'b0;
    end
    else if ( (fsm_output[8]) | (fsm_output[6]) | (fsm_output[4]) | (fsm_output[2])
        | (fsm_output[11]) | (fsm_output[13]) ) begin
      R_21_7_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_3_xor_14_nl, loop_DES_rounds_16_xor_14_cse,
          loop_DES_rounds_7_xor_12_nl, loop_DES_rounds_11_xor_12_cse, loop_DES_rounds_12_xor_14_nl,
          {(fsm_output[2]) , R_or_152_nl , (fsm_output[6]) , (fsm_output[8]) , (fsm_output[11])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_25_6_sva <= 1'b0;
    end
    else if ( (fsm_output[2]) | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[9])
        | (fsm_output[11]) | (fsm_output[13]) ) begin
      R_25_6_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_3_xor_22_nl, loop_DES_rounds_6_xor_20_nl,
          loop_DES_rounds_10_xor_20_cse, loop_DES_rounds_10_xor_22_cse, loop_DES_rounds_16_xor_22_cse,
          {(fsm_output[2]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[9])
          , R_or_133_cse});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_6_5_sva <= 1'b0;
    end
    else if ( (fsm_output[2]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[8])
        ) begin
      R_6_5_sva <= MUX1HOT_s_1_3_2(loop_DES_rounds_3_xor_13_nl, loop_DES_rounds_13_xor_19_cse,
          loop_DES_rounds_11_xor_19_cse, {(fsm_output[2]) , (fsm_output[4]) , R_or_105_cse});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_30_4_sva <= 1'b0;
    end
    else if ( (fsm_output[3]) | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[9])
        | (fsm_output[11]) | (fsm_output[13]) ) begin
      R_30_4_sva <= MUX1HOT_s_1_4_2(loop_DES_rounds_16_xor_30_cse, loop_DES_rounds_10_xor_30_cse,
          loop_DES_rounds_6_xor_19_cse, loop_DES_rounds_16_xor_19_cse, {(fsm_output[3])
          , R_or_cse , (fsm_output[9]) , R_or_133_cse});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_29_4_sva <= 1'b0;
      R_26_4_sva <= 1'b0;
    end
    else if ( R_or_66_cse ) begin
      R_29_4_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_16_xor_28_cse, loop_DES_rounds_10_xor_28_cse,
          loop_DES_rounds_5_xor_21_cse, loop_DES_rounds_15_xor_21_cse, loop_DES_rounds_13_xor_19_cse,
          {(fsm_output[3]) , R_or_cse , (fsm_output[10]) , (fsm_output[12]) , (fsm_output[14])});
      R_26_4_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_4_xor_22_nl, loop_DES_rounds_10_xor_22_cse,
          loop_DES_rounds_7_xor_28_cse, loop_DES_rounds_15_xor_28_cse, loop_DES_rounds_13_xor_30_cse,
          {(fsm_output[3]) , R_or_cse , (fsm_output[10]) , (fsm_output[12]) , (fsm_output[14])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_9_4_sva <= 1'b0;
    end
    else if ( (fsm_output[7]) | (fsm_output[5]) | (fsm_output[3]) ) begin
      R_9_4_sva <= MUX_s_1_2_2(loop_DES_rounds_12_xor_13_cse, loop_DES_rounds_10_xor_13_cse,
          R_or_cse);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      R_22_7_sva <= 1'b0;
    end
    else if ( (fsm_output[3]) | (fsm_output[6]) | (fsm_output[8]) | (fsm_output[10])
        | (fsm_output[12]) | (fsm_output[14]) ) begin
      R_22_7_sva <= MUX1HOT_s_1_5_2(loop_DES_rounds_16_xor_20_cse, loop_DES_rounds_16_xor_14_cse,
          loop_DES_rounds_11_xor_14_cse, loop_DES_rounds_7_xor_22_cse, loop_DES_rounds_13_xor_22_nl,
          {(fsm_output[3]) , (fsm_output[6]) , (fsm_output[8]) , (fsm_output[10])
          , R_or_127_cse});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_input_ftd <= 63'b000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( fsm_output[0] ) begin
      reg_input_ftd <= input_rsci_idat[63:1];
    end
  end
  assign loop_DES_rounds_1_xor_31_nl = (input_rsci_idat[56]) ^ (ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_17[3]);
  assign loop_DES_rounds_2_xor_31_nl = (reg_input_ftd[56]) ^ (s_output_1_3_0_54_sva[3]);
  assign loop_DES_rounds_15_xor_3_nl = R_1_9_sva ^ (O_1_out[0]);
  assign loop_DES_rounds_1_xor_25_nl = (input_rsci_idat[32]) ^ (ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_17[2]);
  assign loop_DES_rounds_2_xor_25_nl = (reg_input_ftd[32]) ^ (s_output_1_3_0_39_sva[2]);
  assign loop_DES_rounds_8_xor_5_nl = R_27_10_sva ^ (O_1_out_7[0]);
  assign loop_DES_rounds_1_xor_11_nl = (input_rsci_idat[42]) ^ (ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_17[1]);
  assign loop_DES_rounds_2_xor_19_nl = (reg_input_ftd[8]) ^ (s_output_1_19_16_5_sva[3]);
  assign loop_DES_rounds_8_xor_11_nl = R_1_9_sva ^ (O_1_out_4[1]);
  assign loop_DES_rounds_12_xor_6_nl = R_1_7_sva ^ (O_1_out_5[2]);
  assign loop_DES_rounds_14_xor_3_nl = R_1_7_sva ^ (O_1_out[0]);
  assign loop_DES_rounds_1_xor_22_nl = (input_rsci_idat[46]) ^ (ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_17[0]);
  assign loop_DES_rounds_2_xor_16_nl = (reg_input_ftd[4]) ^ (s_output_1_19_16_20_sva[3]);
  assign loop_DES_rounds_8_xor_29_nl = R_1_6_sva ^ (O_1_out_3[0]);
  assign loop_DES_rounds_1_xor_17_nl = (input_rsci_idat[0]) ^ (ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_17[1]);
  assign loop_DES_rounds_2_xor_17_nl = (reg_input_ftd[0]) ^ (s_output_1_3_0_24_sva[1]);
  assign loop_DES_rounds_5_xor_3_nl = R_14_3_sva ^ (O_1_out[0]);
  assign loop_DES_rounds_7_xor_6_nl = R_3_1_sva ^ (O_1_out_5[2]);
  assign loop_DES_rounds_1_xor_29_nl = (input_rsci_idat[48]) ^ (O_1_out_3[0]);
  assign loop_DES_rounds_1_xor_2_nl = (input_rsci_idat[60]) ^ (ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_17[2]);
  assign loop_DES_rounds_1_xor_10_nl = (input_rsci_idat[28]) ^ (ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_17[2]);
  assign loop_DES_rounds_2_xor_10_nl = (reg_input_ftd[28]) ^ (s_output_1_3_0_54_sva[2]);
  assign loop_DES_rounds_6_xor_27_nl = R_1_7_sva ^ (O_1_out_6[1]);
  assign loop_DES_rounds_1_xor_4_nl = (input_rsci_idat[52]) ^ (ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_17[1]);
  assign loop_DES_rounds_2_xor_18_nl = (reg_input_ftd[62]) ^ (s_output_1_3_0_24_sva[3]);
  assign loop_DES_rounds_1_xor_6_nl = (input_rsci_idat[44]) ^ (ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_17[2]);
  assign loop_DES_rounds_2_xor_26_nl = (reg_input_ftd[30]) ^ (s_output_1_3_0_39_sva[3]);
  assign loop_DES_rounds_1_xor_24_nl = (input_rsci_idat[38]) ^ (ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_17[3]);
  assign loop_DES_rounds_2_xor_23_nl = (reg_input_ftd[24]) ^ (s_output_1_19_16_35_sva[2]);
  assign loop_DES_rounds_1_xor_9_nl = (input_rsci_idat[34]) ^ (ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_17[0]);
  assign loop_DES_rounds_2_xor_9_nl = (reg_input_ftd[34]) ^ (s_output_1_3_0_9_sva[0]);
  assign loop_DES_rounds_4_xor_14_nl = R_1_7_sva ^ (O_1_out_1[1]);
  assign loop_DES_rounds_7_xor_27_nl = R_10_1_sva ^ (O_1_out_6[1]);
  assign loop_DES_rounds_1_xor_1_nl = (input_rsci_idat[2]) ^ (O_1_out_3[2]);
  assign loop_DES_rounds_2_xor_1_nl = (reg_input_ftd[2]) ^ (s_output_1_19_16_20_sva[2]);
  assign loop_DES_rounds_6_xor_14_nl = R_11_1_sva ^ (O_1_out_1[1]);
  assign loop_DES_rounds_13_xor_20_nl = R_15_1_sva ^ (O_1_out_4[0]);
  assign loop_DES_rounds_1_xor_5_nl = (input_rsci_idat[18]) ^ (ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_17[0]);
  assign loop_DES_rounds_3_xor_7_nl = R_11_3_sva ^ (O_1_out_1[2]);
  assign loop_DES_rounds_13_xor_9_nl = R_11_11_sva ^ (O_1_out_8[0]);
  assign loop_DES_rounds_1_xor_27_nl = (input_rsci_idat[40]) ^ (ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_17[1]);
  assign loop_DES_rounds_3_xor_8_nl = R_16_3_sva ^ (O_1_out[3]);
  assign loop_DES_rounds_5_xor_8_nl = R_19_11_sva ^ (O_1_out[3]);
  assign loop_DES_rounds_1_xor_12_nl = (input_rsci_idat[20]) ^ (ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_17[1]);
  assign loop_DES_rounds_5_xor_10_nl = R_20_11_sva ^ (O_1_out_4[2]);
  assign loop_DES_rounds_1_xor_18_nl = (input_rsci_idat[62]) ^ (ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_17[3]);
  assign loop_DES_rounds_3_xor_16_nl = R_15_9_sva ^ (O_1_out_3[3]);
  assign loop_DES_rounds_5_xor_16_nl = R_23_11_sva ^ (O_1_out_3[3]);
  assign loop_DES_rounds_1_xor_20_nl = (input_rsci_idat[54]) ^ (ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_17[0]);
  assign loop_DES_rounds_3_xor_18_nl = R_23_11_sva ^ (O_1_out_5[3]);
  assign loop_DES_rounds_11_xor_5_nl = R_0_11_sva ^ (O_1_out_7[0]);
  assign loop_DES_rounds_13_xor_6_nl = R_3_3_sva ^ (O_1_out_5[2]);
  assign loop_DES_rounds_1_xor_26_nl = (input_rsci_idat[30]) ^ (ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_17[3]);
  assign loop_DES_rounds_3_xor_24_nl = R_31_4_sva ^ (O_1_out_8[3]);
  assign loop_DES_rounds_5_xor_24_nl = R_27_11_sva ^ (O_1_out_8[3]);
  assign loop_DES_rounds_1_xor_28_nl = (input_rsci_idat[22]) ^ (ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_17[0]);
  assign loop_DES_rounds_3_xor_26_nl = R_27_11_sva ^ (O_1_out_7[3]);
  assign loop_DES_rounds_5_xor_26_nl = R_28_11_sva ^ (O_1_out_7[3]);
  assign loop_DES_rounds_1_xor_21_nl = (input_rsci_idat[16]) ^ (ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_17[2]);
  assign loop_DES_rounds_3_xor_23_nl = R_31_3_sva ^ (O_1_out[2]);
  assign loop_DES_rounds_13_xor_32_nl = R_31_11_sva ^ (O_1_out_1[0]);
  assign loop_DES_rounds_1_xor_13_nl = (input_rsci_idat[50]) ^ (O_1_out_3[1]);
  assign loop_DES_rounds_13_xor_17_nl = R_7_11_sva ^ (O_1_out_5[1]);
  assign loop_DES_rounds_1_xor_15_nl = (input_rsci_idat[58]) ^ (ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_17[3]);
  assign loop_DES_rounds_1_xor_16_nl = (input_rsci_idat[4]) ^ (O_1_out_3[3]);
  assign loop_DES_rounds_13_xor_2_nl = R_15_9_sva ^ (O_1_out_6[2]);
  assign loop_DES_rounds_1_xor_3_nl = (reg_input_ftd[9]) ^ (ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_17[0]);
  assign loop_DES_rounds_3_xor_29_nl = R_0_10_sva ^ (O_1_out_3[0]);
  assign loop_DES_rounds_7_xor_11_nl = R_1_8_sva ^ (O_1_out_4[1]);
  assign loop_DES_rounds_11_xor_31_nl = R_0_9_sva ^ (O_1_out_4[3]);
  assign loop_DES_rounds_13_xor_31_nl = R_0_11_sva ^ (O_1_out_4[3]);
  assign loop_DES_rounds_1_xor_7_nl = (reg_input_ftd[25]) ^ (s_output_1_19_16_20_sva[2]);
  assign loop_DES_rounds_15_xor_5_nl = R_3_3_sva ^ (O_1_out_7[0]);
  assign loop_DES_rounds_1_xor_8_nl = (reg_input_ftd[35]) ^ (ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_17[3]);
  assign loop_DES_rounds_3_xor_2_nl = R_15_10_sva ^ (O_1_out_6[2]);
  assign loop_DES_rounds_1_xor_30_nl = (reg_input_ftd[13]) ^ (ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_17[1]);
  assign loop_DES_rounds_13_xor_5_nl = R_24_3_sva ^ (O_1_out_7[0]);
  assign loop_DES_rounds_1_xor_23_nl = (reg_input_ftd[23]) ^ (ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_17[2]);
  assign loop_DES_rounds_3_xor_32_nl = R_10_10_sva ^ (O_1_out_1[0]);
  assign loop_DES_rounds_11_xor_3_nl = R_12_11_sva ^ (O_1_out[0]);
  assign loop_DES_rounds_14_xor_6_nl = R_10_1_sva ^ (O_1_out_5[2]);
  assign loop_DES_rounds_1_xor_19_nl = (reg_input_ftd[7]) ^ (s_output_1_19_16_20_sva[3]);
  assign loop_DES_rounds_2_xor_6_nl = (reg_input_ftd[44]) ^ (s_output_1_3_0_24_sva[2]);
  assign loop_DES_rounds_6_xor_3_nl = R_31_10_sva ^ (O_1_out[0]);
  assign loop_DES_rounds_9_xor_11_nl = R_0_11_sva ^ (O_1_out_4[1]);
  assign loop_DES_rounds_15_xor_6_nl = R_24_3_sva ^ (O_1_out_5[2]);
  assign R_or_125_nl = (fsm_output[10]) | (fsm_output[12]);
  assign loop_DES_rounds_1_xor_14_nl = (reg_input_ftd[11]) ^ (s_output_1_19_16_20_sva[1]);
  assign loop_DES_rounds_2_xor_8_nl = (reg_input_ftd[36]) ^ (s_output_1_19_16_35_sva[3]);
  assign loop_DES_rounds_4_xor_11_nl = R_0_9_sva ^ (O_1_out_4[1]);
  assign loop_DES_rounds_6_xor_29_nl = R_1_4_sva ^ (O_1_out_3[0]);
  assign loop_DES_rounds_8_xor_3_nl = R_1_4_sva ^ (O_1_out[0]);
  assign loop_DES_rounds_1_xor_32_nl = (reg_input_ftd[5]) ^ (s_output_1_19_16_20_sva[0]);
  assign loop_DES_rounds_3_xor_11_nl = R_10_1_sva ^ (O_1_out_4[1]);
  assign loop_DES_rounds_7_xor_3_nl = R_7_1_sva ^ (O_1_out[0]);
  assign loop_DES_rounds_13_xor_27_nl = R_1_9_sva ^ (O_1_out_6[1]);
  assign R_or_102_nl = (fsm_output[2]) | (fsm_output[9]);
  assign loop_DES_rounds_3_xor_27_nl = R_19_11_sva ^ (O_1_out_6[1]);
  assign loop_DES_rounds_9_xor_27_nl = R_11_1_sva ^ (O_1_out_6[1]);
  assign loop_DES_rounds_13_xor_12_nl = R_2_3_sva ^ (O_1_out_7[1]);
  assign loop_DES_rounds_2_xor_11_nl = (reg_input_ftd[42]) ^ (s_output_1_3_0_54_sva[1]);
  assign loop_DES_rounds_11_xor_29_nl = R_1_9_sva ^ (O_1_out_3[0]);
  assign loop_DES_rounds_3_xor_12_nl = R_20_11_sva ^ (O_1_out_7[1]);
  assign loop_DES_rounds_6_xor_12_nl = R_1_9_sva ^ (O_1_out_7[1]);
  assign loop_DES_rounds_13_xor_14_nl = R_21_3_sva ^ (O_1_out_1[1]);
  assign loop_DES_rounds_3_xor_6_nl = R_27_4_sva ^ (O_1_out_5[2]);
  assign loop_DES_rounds_9_xor_6_nl = R_7_1_sva ^ (O_1_out_5[2]);
  assign loop_DES_rounds_15_xor_27_nl = R_10_10_sva ^ (O_1_out_6[1]);
  assign loop_DES_rounds_3_xor_3_nl = R_0_11_sva ^ (O_1_out[0]);
  assign loop_DES_rounds_5_xor_13_nl = R_6_5_sva ^ (O_1_out_3[1]);
  assign loop_DES_rounds_2_xor_29_nl = (reg_input_ftd[48]) ^ (s_output_1_19_16_20_sva[0]);
  assign loop_DES_rounds_10_xor_29_nl = R_1_8_sva ^ (O_1_out_3[0]);
  assign loop_DES_rounds_2_xor_7_nl = (reg_input_ftd[26]) ^ (s_output_1_19_16_5_sva[2]);
  assign loop_DES_rounds_2_xor_5_nl = (reg_input_ftd[18]) ^ (s_output_1_3_0_39_sva[0]);
  assign loop_DES_rounds_10_xor_5_nl = R_3_1_sva ^ (O_1_out_7[0]);
  assign loop_DES_rounds_2_xor_2_nl = (reg_input_ftd[60]) ^ (s_output_1_19_16_50_sva[2]);
  assign loop_DES_rounds_2_xor_4_nl = (reg_input_ftd[52]) ^ (s_output_1_3_0_9_sva[1]);
  assign loop_DES_rounds_10_xor_4_nl = R_20_1_sva ^ (O_1_out_8[1]);
  assign loop_DES_rounds_2_xor_27_nl = (reg_input_ftd[40]) ^ (s_output_1_19_16_50_sva[1]);
  assign loop_DES_rounds_10_xor_27_nl = R_31_10_sva ^ (O_1_out_6[1]);
  assign loop_DES_rounds_2_xor_12_nl = (reg_input_ftd[20]) ^ (s_output_1_3_0_39_sva[1]);
  assign loop_DES_rounds_2_xor_20_nl = (reg_input_ftd[54]) ^ (s_output_1_3_0_54_sva[0]);
  assign loop_DES_rounds_2_xor_24_nl = (reg_input_ftd[38]) ^ (s_output_1_3_0_9_sva[3]);
  assign loop_DES_rounds_4_xor_6_nl = R_1_4_sva ^ (O_1_out_5[2]);
  assign loop_DES_rounds_6_xor_5_nl = R_20_1_sva ^ (O_1_out_7[0]);
  assign loop_DES_rounds_8_xor_6_nl = R_31_10_sva ^ (O_1_out_5[2]);
  assign loop_DES_rounds_2_xor_28_nl = (reg_input_ftd[22]) ^ (s_output_1_3_0_24_sva[0]);
  assign loop_DES_rounds_2_xor_30_nl = (reg_input_ftd[14]) ^ (s_output_1_19_16_35_sva[1]);
  assign loop_DES_rounds_2_xor_32_nl = (reg_input_ftd[6]) ^ (s_output_1_19_16_5_sva[0]);
  assign loop_DES_rounds_8_xor_27_nl = R_20_1_sva ^ (O_1_out_6[1]);
  assign loop_DES_rounds_2_xor_21_nl = (reg_input_ftd[16]) ^ (s_output_1_3_0_9_sva[2]);
  assign loop_DES_rounds_2_xor_15_nl = (reg_input_ftd[58]) ^ (s_output_1_19_16_50_sva[3]);
  assign loop_DES_rounds_2_xor_13_nl = (reg_input_ftd[50]) ^ (s_output_1_19_16_20_sva[1]);
  assign loop_DES_rounds_2_xor_3_nl = (reg_input_ftd[10]) ^ (s_output_1_19_16_35_sva[0]);
  assign loop_DES_rounds_4_xor_19_nl = R_10_1_sva ^ (O_1_out_1[3]);
  assign loop_DES_rounds_10_xor_3_nl = R_1_6_sva ^ (O_1_out[0]);
  assign loop_DES_rounds_3_xor_5_nl = R_11_11_sva ^ (O_1_out_7[0]);
  assign loop_DES_rounds_9_xor_3_nl = R_10_10_sva ^ (O_1_out[0]);
  assign loop_DES_rounds_13_xor_7_nl = R_12_11_sva ^ (O_1_out_1[2]);
  assign R_or_99_nl = (fsm_output[4]) | (fsm_output[6]);
  assign loop_DES_rounds_3_xor_4_nl = R_23_4_sva ^ (O_1_out_8[1]);
  assign loop_DES_rounds_11_xor_1_nl = R_15_9_sva ^ (O_1_out_3[2]);
  assign loop_DES_rounds_13_xor_1_nl = R_15_11_sva ^ (O_1_out_3[2]);
  assign loop_DES_rounds_3_xor_20_nl = R_24_3_sva ^ (O_1_out_4[0]);
  assign loop_DES_rounds_13_xor_18_nl = R_24_11_sva ^ (O_1_out_5[3]);
  assign loop_DES_rounds_3_xor_30_nl = R_3_3_sva ^ (O_1_out[1]);
  assign loop_DES_rounds_13_xor_25_nl = R_3_11_sva ^ (O_1_out_7[2]);
  assign loop_DES_rounds_3_xor_21_nl = R_31_11_sva ^ (O_1_out_8[2]);
  assign loop_DES_rounds_13_xor_23_nl = R_4_11_sva ^ (O_1_out[2]);
  assign loop_DES_rounds_3_xor_28_nl = R_28_11_sva ^ (O_1_out_5[0]);
  assign loop_DES_rounds_3_xor_19_nl = R_1_4_sva ^ (O_1_out_1[3]);
  assign loop_DES_rounds_5_xor_28_nl = R_26_5_sva ^ (O_1_out_5[0]);
  assign loop_DES_rounds_2_xor_14_nl = (reg_input_ftd[12]) ^ (s_output_1_19_16_5_sva[1]);
  assign loop_DES_rounds_14_xor_11_nl = R_1_14_sva ^ (O_1_out_4[1]);
  assign loop_DES_rounds_2_xor_22_nl = (reg_input_ftd[46]) ^ (s_output_1_19_16_50_sva[0]);
  assign loop_DES_rounds_6_xor_11_nl = R_1_6_sva ^ (O_1_out_4[1]);
  assign loop_DES_rounds_9_xor_29_nl = R_1_7_sva ^ (O_1_out_3[0]);
  assign loop_DES_rounds_13_xor_3_nl = R_31_3_sva ^ (O_1_out[0]);
  assign loop_DES_rounds_3_xor_14_nl = R_1_6_sva ^ (O_1_out_1[1]);
  assign loop_DES_rounds_7_xor_12_nl = R_10_10_sva ^ (O_1_out_7[1]);
  assign loop_DES_rounds_12_xor_14_nl = R_10_1_sva ^ (O_1_out_1[1]);
  assign R_or_152_nl = (fsm_output[4]) | (fsm_output[13]);
  assign loop_DES_rounds_3_xor_22_nl = R_1_8_sva ^ (O_1_out_6[0]);
  assign loop_DES_rounds_6_xor_20_nl = R_22_7_sva ^ (O_1_out_4[0]);
  assign loop_DES_rounds_3_xor_13_nl = R_7_11_sva ^ (O_1_out_3[1]);
  assign loop_DES_rounds_4_xor_22_nl = R_1_9_sva ^ (O_1_out_6[0]);
  assign loop_DES_rounds_13_xor_22_nl = R_22_7_sva ^ (O_1_out_6[0]);

  function automatic [0:0] MUX1HOT_s_1_14_2;
    input [0:0] input_13;
    input [0:0] input_12;
    input [0:0] input_11;
    input [0:0] input_10;
    input [0:0] input_9;
    input [0:0] input_8;
    input [0:0] input_7;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [13:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    result = result | ( input_7 & {1{sel[7]}});
    result = result | ( input_8 & {1{sel[8]}});
    result = result | ( input_9 & {1{sel[9]}});
    result = result | ( input_10 & {1{sel[10]}});
    result = result | ( input_11 & {1{sel[11]}});
    result = result | ( input_12 & {1{sel[12]}});
    result = result | ( input_13 & {1{sel[13]}});
    MUX1HOT_s_1_14_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_15_2;
    input [0:0] input_14;
    input [0:0] input_13;
    input [0:0] input_12;
    input [0:0] input_11;
    input [0:0] input_10;
    input [0:0] input_9;
    input [0:0] input_8;
    input [0:0] input_7;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [14:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    result = result | ( input_7 & {1{sel[7]}});
    result = result | ( input_8 & {1{sel[8]}});
    result = result | ( input_9 & {1{sel[9]}});
    result = result | ( input_10 & {1{sel[10]}});
    result = result | ( input_11 & {1{sel[11]}});
    result = result | ( input_12 & {1{sel[12]}});
    result = result | ( input_13 & {1{sel[13]}});
    result = result | ( input_14 & {1{sel[14]}});
    MUX1HOT_s_1_15_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_5_2;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [4:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_6_2;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [5:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    MUX1HOT_s_1_6_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_7_2;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [6:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    des_check
// ------------------------------------------------------------------


module des_check (
  clk, rst, input_rsc_dat, input_rsc_triosy_lz, key_rsc_dat, key_rsc_triosy_lz, return_rsc_dat,
      return_rsc_triosy_lz
);
  input clk;
  input rst;
  input [63:0] input_rsc_dat;
  output input_rsc_triosy_lz;
  input [63:0] key_rsc_dat;
  output key_rsc_triosy_lz;
  output [63:0] return_rsc_dat;
  output return_rsc_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  des_check_core des_check_core_inst (
      .clk(clk),
      .rst(rst),
      .input_rsc_dat(input_rsc_dat),
      .input_rsc_triosy_lz(input_rsc_triosy_lz),
      .key_rsc_dat(key_rsc_dat),
      .key_rsc_triosy_lz(key_rsc_triosy_lz),
      .return_rsc_dat(return_rsc_dat),
      .return_rsc_triosy_lz(return_rsc_triosy_lz)
    );
endmodule



