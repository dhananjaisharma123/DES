
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ../td_ccore_solutions/ROM_1i6_1o4_ef4da7ff735c86ba85f23e51741d972cb3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Mon Mar  1 00:26:55 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i6_1o4_ef4da7ff735c86ba85f23e51741d972cb3
// ------------------------------------------------------------------


module ROM_1i6_1o4_ef4da7ff735c86ba85f23e51741d972cb3 (
  I_1, O_1
);
  input [5:0] I_1;
  output [3:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_4_64_2(4'b1101, 4'b0010, 4'b1000, 4'b0100, 4'b0110, 4'b1111,
      4'b1011, 4'b0001, 4'b1010, 4'b1001, 4'b0011, 4'b1110, 4'b0101, 4'b0000, 4'b1100,
      4'b0111, 4'b0001, 4'b1111, 4'b1101, 4'b1000, 4'b1010, 4'b0011, 4'b0111, 4'b0100,
      4'b1100, 4'b0101, 4'b0110, 4'b1011, 4'b0000, 4'b1110, 4'b1001, 4'b0010, 4'b0111,
      4'b1011, 4'b0100, 4'b0001, 4'b1001, 4'b1100, 4'b1110, 4'b0010, 4'b0000, 4'b0110,
      4'b1010, 4'b1101, 4'b1111, 4'b0011, 4'b0101, 4'b1000, 4'b0010, 4'b0001, 4'b1110,
      4'b0111, 4'b0100, 4'b1010, 4'b1000, 4'b1101, 4'b1111, 4'b1100, 4'b1001, 4'b0000,
      4'b0011, 4'b0101, 4'b0110, 4'b1011, I_1);

  function automatic [3:0] MUX_v_4_64_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [3:0] input_8;
    input [3:0] input_9;
    input [3:0] input_10;
    input [3:0] input_11;
    input [3:0] input_12;
    input [3:0] input_13;
    input [3:0] input_14;
    input [3:0] input_15;
    input [3:0] input_16;
    input [3:0] input_17;
    input [3:0] input_18;
    input [3:0] input_19;
    input [3:0] input_20;
    input [3:0] input_21;
    input [3:0] input_22;
    input [3:0] input_23;
    input [3:0] input_24;
    input [3:0] input_25;
    input [3:0] input_26;
    input [3:0] input_27;
    input [3:0] input_28;
    input [3:0] input_29;
    input [3:0] input_30;
    input [3:0] input_31;
    input [3:0] input_32;
    input [3:0] input_33;
    input [3:0] input_34;
    input [3:0] input_35;
    input [3:0] input_36;
    input [3:0] input_37;
    input [3:0] input_38;
    input [3:0] input_39;
    input [3:0] input_40;
    input [3:0] input_41;
    input [3:0] input_42;
    input [3:0] input_43;
    input [3:0] input_44;
    input [3:0] input_45;
    input [3:0] input_46;
    input [3:0] input_47;
    input [3:0] input_48;
    input [3:0] input_49;
    input [3:0] input_50;
    input [3:0] input_51;
    input [3:0] input_52;
    input [3:0] input_53;
    input [3:0] input_54;
    input [3:0] input_55;
    input [3:0] input_56;
    input [3:0] input_57;
    input [3:0] input_58;
    input [3:0] input_59;
    input [3:0] input_60;
    input [3:0] input_61;
    input [3:0] input_62;
    input [3:0] input_63;
    input [5:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_4_64_2 = result;
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i6_1o4_d0e242163cbb0b2ce9c4399bc1cb50f5b3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Mon Mar  1 00:26:47 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i6_1o4_d0e242163cbb0b2ce9c4399bc1cb50f5b3
// ------------------------------------------------------------------


module ROM_1i6_1o4_d0e242163cbb0b2ce9c4399bc1cb50f5b3 (
  I_1, O_1
);
  input [5:0] I_1;
  output [3:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_4_64_2(4'b0111, 4'b1101, 4'b1110, 4'b0011, 4'b0000, 4'b0110,
      4'b1001, 4'b1010, 4'b0001, 4'b0010, 4'b1000, 4'b0101, 4'b1011, 4'b1100, 4'b0100,
      4'b1111, 4'b1101, 4'b1000, 4'b1011, 4'b0101, 4'b0110, 4'b1111, 4'b0000, 4'b0011,
      4'b0100, 4'b0111, 4'b0010, 4'b1100, 4'b0001, 4'b1010, 4'b1110, 4'b1001, 4'b1010,
      4'b0110, 4'b1001, 4'b0000, 4'b1100, 4'b1011, 4'b0111, 4'b1101, 4'b1111, 4'b0001,
      4'b0011, 4'b1110, 4'b0101, 4'b0010, 4'b1000, 4'b0100, 4'b0011, 4'b1111, 4'b0000,
      4'b0110, 4'b1010, 4'b0001, 4'b1101, 4'b1000, 4'b1001, 4'b0100, 4'b0101, 4'b1011,
      4'b1100, 4'b0111, 4'b0010, 4'b1110, I_1);

  function automatic [3:0] MUX_v_4_64_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [3:0] input_8;
    input [3:0] input_9;
    input [3:0] input_10;
    input [3:0] input_11;
    input [3:0] input_12;
    input [3:0] input_13;
    input [3:0] input_14;
    input [3:0] input_15;
    input [3:0] input_16;
    input [3:0] input_17;
    input [3:0] input_18;
    input [3:0] input_19;
    input [3:0] input_20;
    input [3:0] input_21;
    input [3:0] input_22;
    input [3:0] input_23;
    input [3:0] input_24;
    input [3:0] input_25;
    input [3:0] input_26;
    input [3:0] input_27;
    input [3:0] input_28;
    input [3:0] input_29;
    input [3:0] input_30;
    input [3:0] input_31;
    input [3:0] input_32;
    input [3:0] input_33;
    input [3:0] input_34;
    input [3:0] input_35;
    input [3:0] input_36;
    input [3:0] input_37;
    input [3:0] input_38;
    input [3:0] input_39;
    input [3:0] input_40;
    input [3:0] input_41;
    input [3:0] input_42;
    input [3:0] input_43;
    input [3:0] input_44;
    input [3:0] input_45;
    input [3:0] input_46;
    input [3:0] input_47;
    input [3:0] input_48;
    input [3:0] input_49;
    input [3:0] input_50;
    input [3:0] input_51;
    input [3:0] input_52;
    input [3:0] input_53;
    input [3:0] input_54;
    input [3:0] input_55;
    input [3:0] input_56;
    input [3:0] input_57;
    input [3:0] input_58;
    input [3:0] input_59;
    input [3:0] input_60;
    input [3:0] input_61;
    input [3:0] input_62;
    input [3:0] input_63;
    input [5:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_4_64_2 = result;
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i6_1o4_752c7ca65a598ada4acee0cd63d199c3b3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Mon Mar  1 00:26:38 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i6_1o4_752c7ca65a598ada4acee0cd63d199c3b3
// ------------------------------------------------------------------


module ROM_1i6_1o4_752c7ca65a598ada4acee0cd63d199c3b3 (
  I_1, O_1
);
  input [5:0] I_1;
  output [3:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_4_64_2(4'b0100, 4'b1011, 4'b0010, 4'b1110, 4'b1111, 4'b0000,
      4'b1000, 4'b1101, 4'b0011, 4'b1100, 4'b1001, 4'b0111, 4'b0101, 4'b1010, 4'b0110,
      4'b0001, 4'b1101, 4'b0000, 4'b1011, 4'b0111, 4'b0100, 4'b1001, 4'b0001, 4'b1010,
      4'b1110, 4'b0011, 4'b0101, 4'b1100, 4'b0010, 4'b1111, 4'b1000, 4'b0110, 4'b0001,
      4'b0100, 4'b1011, 4'b1101, 4'b1100, 4'b0011, 4'b0111, 4'b1110, 4'b1010, 4'b1111,
      4'b0110, 4'b1000, 4'b0000, 4'b0101, 4'b1001, 4'b0010, 4'b0110, 4'b1011, 4'b1101,
      4'b1000, 4'b0001, 4'b0100, 4'b1010, 4'b0111, 4'b1001, 4'b0101, 4'b0000, 4'b1111,
      4'b1110, 4'b0010, 4'b0011, 4'b1100, I_1);

  function automatic [3:0] MUX_v_4_64_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [3:0] input_8;
    input [3:0] input_9;
    input [3:0] input_10;
    input [3:0] input_11;
    input [3:0] input_12;
    input [3:0] input_13;
    input [3:0] input_14;
    input [3:0] input_15;
    input [3:0] input_16;
    input [3:0] input_17;
    input [3:0] input_18;
    input [3:0] input_19;
    input [3:0] input_20;
    input [3:0] input_21;
    input [3:0] input_22;
    input [3:0] input_23;
    input [3:0] input_24;
    input [3:0] input_25;
    input [3:0] input_26;
    input [3:0] input_27;
    input [3:0] input_28;
    input [3:0] input_29;
    input [3:0] input_30;
    input [3:0] input_31;
    input [3:0] input_32;
    input [3:0] input_33;
    input [3:0] input_34;
    input [3:0] input_35;
    input [3:0] input_36;
    input [3:0] input_37;
    input [3:0] input_38;
    input [3:0] input_39;
    input [3:0] input_40;
    input [3:0] input_41;
    input [3:0] input_42;
    input [3:0] input_43;
    input [3:0] input_44;
    input [3:0] input_45;
    input [3:0] input_46;
    input [3:0] input_47;
    input [3:0] input_48;
    input [3:0] input_49;
    input [3:0] input_50;
    input [3:0] input_51;
    input [3:0] input_52;
    input [3:0] input_53;
    input [3:0] input_54;
    input [3:0] input_55;
    input [3:0] input_56;
    input [3:0] input_57;
    input [3:0] input_58;
    input [3:0] input_59;
    input [3:0] input_60;
    input [3:0] input_61;
    input [3:0] input_62;
    input [3:0] input_63;
    input [5:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_4_64_2 = result;
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i6_1o4_3c5c29b75c561d2b741f22e5a3a569dbb3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Mon Mar  1 00:26:30 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i6_1o4_3c5c29b75c561d2b741f22e5a3a569dbb3
// ------------------------------------------------------------------


module ROM_1i6_1o4_3c5c29b75c561d2b741f22e5a3a569dbb3 (
  I_1, O_1
);
  input [5:0] I_1;
  output [3:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_4_64_2(4'b1010, 4'b0000, 4'b1001, 4'b1110, 4'b0110, 4'b0011,
      4'b1111, 4'b0101, 4'b0001, 4'b1101, 4'b1100, 4'b0111, 4'b1011, 4'b0100, 4'b0010,
      4'b1000, 4'b1101, 4'b0111, 4'b0000, 4'b1001, 4'b0011, 4'b0100, 4'b0110, 4'b1010,
      4'b0010, 4'b1000, 4'b0101, 4'b1110, 4'b1100, 4'b1011, 4'b1111, 4'b0001, 4'b1101,
      4'b0110, 4'b0100, 4'b1001, 4'b1000, 4'b1111, 4'b0011, 4'b0000, 4'b1011, 4'b0001,
      4'b0010, 4'b1100, 4'b0101, 4'b1010, 4'b1110, 4'b0111, 4'b0001, 4'b1010, 4'b1101,
      4'b0000, 4'b0110, 4'b1001, 4'b1000, 4'b0111, 4'b0100, 4'b1111, 4'b1110, 4'b0011,
      4'b1011, 4'b0101, 4'b0010, 4'b1100, I_1);

  function automatic [3:0] MUX_v_4_64_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [3:0] input_8;
    input [3:0] input_9;
    input [3:0] input_10;
    input [3:0] input_11;
    input [3:0] input_12;
    input [3:0] input_13;
    input [3:0] input_14;
    input [3:0] input_15;
    input [3:0] input_16;
    input [3:0] input_17;
    input [3:0] input_18;
    input [3:0] input_19;
    input [3:0] input_20;
    input [3:0] input_21;
    input [3:0] input_22;
    input [3:0] input_23;
    input [3:0] input_24;
    input [3:0] input_25;
    input [3:0] input_26;
    input [3:0] input_27;
    input [3:0] input_28;
    input [3:0] input_29;
    input [3:0] input_30;
    input [3:0] input_31;
    input [3:0] input_32;
    input [3:0] input_33;
    input [3:0] input_34;
    input [3:0] input_35;
    input [3:0] input_36;
    input [3:0] input_37;
    input [3:0] input_38;
    input [3:0] input_39;
    input [3:0] input_40;
    input [3:0] input_41;
    input [3:0] input_42;
    input [3:0] input_43;
    input [3:0] input_44;
    input [3:0] input_45;
    input [3:0] input_46;
    input [3:0] input_47;
    input [3:0] input_48;
    input [3:0] input_49;
    input [3:0] input_50;
    input [3:0] input_51;
    input [3:0] input_52;
    input [3:0] input_53;
    input [3:0] input_54;
    input [3:0] input_55;
    input [3:0] input_56;
    input [3:0] input_57;
    input [3:0] input_58;
    input [3:0] input_59;
    input [3:0] input_60;
    input [3:0] input_61;
    input [3:0] input_62;
    input [3:0] input_63;
    input [5:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_4_64_2 = result;
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i6_1o4_51ba7157b272cd3b87451219caf38e7cb3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Mon Mar  1 00:26:22 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i6_1o4_51ba7157b272cd3b87451219caf38e7cb3
// ------------------------------------------------------------------


module ROM_1i6_1o4_51ba7157b272cd3b87451219caf38e7cb3 (
  I_1, O_1
);
  input [5:0] I_1;
  output [3:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_4_64_2(4'b1100, 4'b0001, 4'b1010, 4'b1111, 4'b1001, 4'b0010,
      4'b0110, 4'b1000, 4'b0000, 4'b1101, 4'b0011, 4'b0100, 4'b1110, 4'b0111, 4'b0101,
      4'b1011, 4'b1010, 4'b1111, 4'b0100, 4'b0010, 4'b0111, 4'b1100, 4'b1001, 4'b0101,
      4'b0110, 4'b0001, 4'b1101, 4'b1110, 4'b0000, 4'b1011, 4'b0011, 4'b1000, 4'b1001,
      4'b1110, 4'b1111, 4'b0101, 4'b0010, 4'b1000, 4'b1100, 4'b0011, 4'b0111, 4'b0000,
      4'b0100, 4'b1010, 4'b0001, 4'b1101, 4'b1011, 4'b0110, 4'b0100, 4'b0011, 4'b0010,
      4'b1100, 4'b1001, 4'b0101, 4'b1111, 4'b1010, 4'b1011, 4'b1110, 4'b0001, 4'b0111,
      4'b0110, 4'b0000, 4'b1000, 4'b1101, I_1);

  function automatic [3:0] MUX_v_4_64_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [3:0] input_8;
    input [3:0] input_9;
    input [3:0] input_10;
    input [3:0] input_11;
    input [3:0] input_12;
    input [3:0] input_13;
    input [3:0] input_14;
    input [3:0] input_15;
    input [3:0] input_16;
    input [3:0] input_17;
    input [3:0] input_18;
    input [3:0] input_19;
    input [3:0] input_20;
    input [3:0] input_21;
    input [3:0] input_22;
    input [3:0] input_23;
    input [3:0] input_24;
    input [3:0] input_25;
    input [3:0] input_26;
    input [3:0] input_27;
    input [3:0] input_28;
    input [3:0] input_29;
    input [3:0] input_30;
    input [3:0] input_31;
    input [3:0] input_32;
    input [3:0] input_33;
    input [3:0] input_34;
    input [3:0] input_35;
    input [3:0] input_36;
    input [3:0] input_37;
    input [3:0] input_38;
    input [3:0] input_39;
    input [3:0] input_40;
    input [3:0] input_41;
    input [3:0] input_42;
    input [3:0] input_43;
    input [3:0] input_44;
    input [3:0] input_45;
    input [3:0] input_46;
    input [3:0] input_47;
    input [3:0] input_48;
    input [3:0] input_49;
    input [3:0] input_50;
    input [3:0] input_51;
    input [3:0] input_52;
    input [3:0] input_53;
    input [3:0] input_54;
    input [3:0] input_55;
    input [3:0] input_56;
    input [3:0] input_57;
    input [3:0] input_58;
    input [3:0] input_59;
    input [3:0] input_60;
    input [3:0] input_61;
    input [3:0] input_62;
    input [3:0] input_63;
    input [5:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_4_64_2 = result;
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i6_1o4_cfafff97e973ca9580e646fecdc2f814b3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Mon Mar  1 00:26:13 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i6_1o4_cfafff97e973ca9580e646fecdc2f814b3
// ------------------------------------------------------------------


module ROM_1i6_1o4_cfafff97e973ca9580e646fecdc2f814b3 (
  I_1, O_1
);
  input [5:0] I_1;
  output [3:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_4_64_2(4'b1111, 4'b0001, 4'b1000, 4'b1110, 4'b0110, 4'b1011,
      4'b0011, 4'b0100, 4'b1001, 4'b0111, 4'b0010, 4'b1101, 4'b1100, 4'b0000, 4'b0101,
      4'b1010, 4'b0011, 4'b1101, 4'b0100, 4'b0111, 4'b1111, 4'b0010, 4'b1000, 4'b1110,
      4'b1100, 4'b0000, 4'b0001, 4'b1010, 4'b0110, 4'b1001, 4'b1011, 4'b0101, 4'b0000,
      4'b1110, 4'b0111, 4'b1011, 4'b1010, 4'b0100, 4'b1101, 4'b0001, 4'b0101, 4'b1000,
      4'b1100, 4'b0110, 4'b1001, 4'b0011, 4'b0010, 4'b1111, 4'b1101, 4'b1000, 4'b1010,
      4'b0001, 4'b0011, 4'b1111, 4'b0100, 4'b0010, 4'b1011, 4'b0110, 4'b0111, 4'b1100,
      4'b0000, 4'b0101, 4'b1110, 4'b1001, I_1);

  function automatic [3:0] MUX_v_4_64_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [3:0] input_8;
    input [3:0] input_9;
    input [3:0] input_10;
    input [3:0] input_11;
    input [3:0] input_12;
    input [3:0] input_13;
    input [3:0] input_14;
    input [3:0] input_15;
    input [3:0] input_16;
    input [3:0] input_17;
    input [3:0] input_18;
    input [3:0] input_19;
    input [3:0] input_20;
    input [3:0] input_21;
    input [3:0] input_22;
    input [3:0] input_23;
    input [3:0] input_24;
    input [3:0] input_25;
    input [3:0] input_26;
    input [3:0] input_27;
    input [3:0] input_28;
    input [3:0] input_29;
    input [3:0] input_30;
    input [3:0] input_31;
    input [3:0] input_32;
    input [3:0] input_33;
    input [3:0] input_34;
    input [3:0] input_35;
    input [3:0] input_36;
    input [3:0] input_37;
    input [3:0] input_38;
    input [3:0] input_39;
    input [3:0] input_40;
    input [3:0] input_41;
    input [3:0] input_42;
    input [3:0] input_43;
    input [3:0] input_44;
    input [3:0] input_45;
    input [3:0] input_46;
    input [3:0] input_47;
    input [3:0] input_48;
    input [3:0] input_49;
    input [3:0] input_50;
    input [3:0] input_51;
    input [3:0] input_52;
    input [3:0] input_53;
    input [3:0] input_54;
    input [3:0] input_55;
    input [3:0] input_56;
    input [3:0] input_57;
    input [3:0] input_58;
    input [3:0] input_59;
    input [3:0] input_60;
    input [3:0] input_61;
    input [3:0] input_62;
    input [3:0] input_63;
    input [5:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_4_64_2 = result;
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i6_1o4_ef717c7c87dc90ac6f7b34d533fe115fb3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Mon Mar  1 00:26:05 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i6_1o4_ef717c7c87dc90ac6f7b34d533fe115fb3
// ------------------------------------------------------------------


module ROM_1i6_1o4_ef717c7c87dc90ac6f7b34d533fe115fb3 (
  I_1, O_1
);
  input [5:0] I_1;
  output [3:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_4_64_2(4'b0010, 4'b1100, 4'b0100, 4'b0001, 4'b0111, 4'b1010,
      4'b1011, 4'b0110, 4'b1000, 4'b0101, 4'b0011, 4'b1111, 4'b1101, 4'b0000, 4'b1110,
      4'b1001, 4'b1110, 4'b1011, 4'b0010, 4'b1100, 4'b0100, 4'b0111, 4'b1101, 4'b0001,
      4'b0101, 4'b0000, 4'b1111, 4'b1010, 4'b0011, 4'b1001, 4'b1000, 4'b0110, 4'b0100,
      4'b0010, 4'b0001, 4'b1011, 4'b1010, 4'b1101, 4'b0111, 4'b1000, 4'b1111, 4'b1001,
      4'b1100, 4'b0101, 4'b0110, 4'b0011, 4'b0000, 4'b1110, 4'b1011, 4'b1000, 4'b1100,
      4'b0111, 4'b0001, 4'b1110, 4'b0010, 4'b1101, 4'b0110, 4'b1111, 4'b0000, 4'b1001,
      4'b1010, 4'b0100, 4'b0101, 4'b0011, I_1);

  function automatic [3:0] MUX_v_4_64_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [3:0] input_8;
    input [3:0] input_9;
    input [3:0] input_10;
    input [3:0] input_11;
    input [3:0] input_12;
    input [3:0] input_13;
    input [3:0] input_14;
    input [3:0] input_15;
    input [3:0] input_16;
    input [3:0] input_17;
    input [3:0] input_18;
    input [3:0] input_19;
    input [3:0] input_20;
    input [3:0] input_21;
    input [3:0] input_22;
    input [3:0] input_23;
    input [3:0] input_24;
    input [3:0] input_25;
    input [3:0] input_26;
    input [3:0] input_27;
    input [3:0] input_28;
    input [3:0] input_29;
    input [3:0] input_30;
    input [3:0] input_31;
    input [3:0] input_32;
    input [3:0] input_33;
    input [3:0] input_34;
    input [3:0] input_35;
    input [3:0] input_36;
    input [3:0] input_37;
    input [3:0] input_38;
    input [3:0] input_39;
    input [3:0] input_40;
    input [3:0] input_41;
    input [3:0] input_42;
    input [3:0] input_43;
    input [3:0] input_44;
    input [3:0] input_45;
    input [3:0] input_46;
    input [3:0] input_47;
    input [3:0] input_48;
    input [3:0] input_49;
    input [3:0] input_50;
    input [3:0] input_51;
    input [3:0] input_52;
    input [3:0] input_53;
    input [3:0] input_54;
    input [3:0] input_55;
    input [3:0] input_56;
    input [3:0] input_57;
    input [3:0] input_58;
    input [3:0] input_59;
    input [3:0] input_60;
    input [3:0] input_61;
    input [3:0] input_62;
    input [3:0] input_63;
    input [5:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_4_64_2 = result;
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i6_1o4_8f60b2fc4a3ee4cef30040071bc0219cb3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Mon Mar  1 00:25:55 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i6_1o4_8f60b2fc4a3ee4cef30040071bc0219cb3
// ------------------------------------------------------------------


module ROM_1i6_1o4_8f60b2fc4a3ee4cef30040071bc0219cb3 (
  I_1, O_1
);
  input [5:0] I_1;
  output [3:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_4_64_2(4'b1110, 4'b0100, 4'b1101, 4'b0001, 4'b0010, 4'b1111,
      4'b1011, 4'b1000, 4'b0011, 4'b1010, 4'b0110, 4'b1100, 4'b0101, 4'b1001, 4'b0000,
      4'b0111, 4'b0000, 4'b1111, 4'b0111, 4'b0100, 4'b1110, 4'b0010, 4'b1101, 4'b0001,
      4'b1010, 4'b0110, 4'b1100, 4'b1011, 4'b1001, 4'b0101, 4'b0011, 4'b1000, 4'b0100,
      4'b0001, 4'b1110, 4'b1000, 4'b1101, 4'b0110, 4'b0010, 4'b1011, 4'b1111, 4'b1100,
      4'b1001, 4'b0111, 4'b0011, 4'b1010, 4'b0101, 4'b0000, 4'b1111, 4'b1100, 4'b1000,
      4'b0010, 4'b0100, 4'b1001, 4'b0001, 4'b0111, 4'b0101, 4'b1011, 4'b0011, 4'b1110,
      4'b1010, 4'b0000, 4'b0110, 4'b1101, I_1);

  function automatic [3:0] MUX_v_4_64_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [3:0] input_8;
    input [3:0] input_9;
    input [3:0] input_10;
    input [3:0] input_11;
    input [3:0] input_12;
    input [3:0] input_13;
    input [3:0] input_14;
    input [3:0] input_15;
    input [3:0] input_16;
    input [3:0] input_17;
    input [3:0] input_18;
    input [3:0] input_19;
    input [3:0] input_20;
    input [3:0] input_21;
    input [3:0] input_22;
    input [3:0] input_23;
    input [3:0] input_24;
    input [3:0] input_25;
    input [3:0] input_26;
    input [3:0] input_27;
    input [3:0] input_28;
    input [3:0] input_29;
    input [3:0] input_30;
    input [3:0] input_31;
    input [3:0] input_32;
    input [3:0] input_33;
    input [3:0] input_34;
    input [3:0] input_35;
    input [3:0] input_36;
    input [3:0] input_37;
    input [3:0] input_38;
    input [3:0] input_39;
    input [3:0] input_40;
    input [3:0] input_41;
    input [3:0] input_42;
    input [3:0] input_43;
    input [3:0] input_44;
    input [3:0] input_45;
    input [3:0] input_46;
    input [3:0] input_47;
    input [3:0] input_48;
    input [3:0] input_49;
    input [3:0] input_50;
    input [3:0] input_51;
    input [3:0] input_52;
    input [3:0] input_53;
    input [3:0] input_54;
    input [3:0] input_55;
    input [3:0] input_56;
    input [3:0] input_57;
    input [3:0] input_58;
    input [3:0] input_59;
    input [3:0] input_60;
    input [3:0] input_61;
    input [3:0] input_62;
    input [3:0] input_63;
    input [5:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_4_64_2 = result;
  end
  endfunction

endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ds6365@hansolo.poly.edu
//  Generated date: Sun Mar 21 13:03:40 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    des_check_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module des_check_core_core_fsm (
  clk, rst, fsm_output, loop_DES_rounds_C_0_tr0
);
  input clk;
  input rst;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;
  input loop_DES_rounds_C_0_tr0;


  // FSM State Type Declaration for des_check_core_core_fsm_1
  parameter
    main_C_0 = 2'd0,
    loop_DES_rounds_C_0 = 2'd1,
    main_C_1 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : des_check_core_core_fsm_1
    case (state_var)
      loop_DES_rounds_C_0 : begin
        fsm_output = 3'b010;
        if ( loop_DES_rounds_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = loop_DES_rounds_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 3'b100;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 3'b001;
        state_var_NS = loop_DES_rounds_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    des_check_core
// ------------------------------------------------------------------


module des_check_core (
  clk, rst, input_rsc_dat, input_rsc_triosy_lz, key_rsc_dat, key_rsc_triosy_lz, return_rsc_dat,
      return_rsc_triosy_lz
);
  input clk;
  input rst;
  input [63:0] input_rsc_dat;
  output input_rsc_triosy_lz;
  input [63:0] key_rsc_dat;
  output key_rsc_triosy_lz;
  output [63:0] return_rsc_dat;
  output return_rsc_triosy_lz;


  // Interconnect Declarations
  wire [63:0] input_rsci_idat;
  wire [63:0] key_rsci_idat;
  reg return_rsci_idat_63;
  reg return_rsci_idat_62;
  reg return_rsci_idat_61;
  reg return_rsci_idat_60;
  reg return_rsci_idat_59;
  reg return_rsci_idat_58;
  reg return_rsci_idat_57;
  reg return_rsci_idat_56;
  reg return_rsci_idat_55;
  reg return_rsci_idat_54;
  reg return_rsci_idat_53;
  reg return_rsci_idat_52;
  reg return_rsci_idat_51;
  reg return_rsci_idat_50;
  reg return_rsci_idat_49;
  reg return_rsci_idat_48;
  reg return_rsci_idat_47;
  reg return_rsci_idat_46;
  reg return_rsci_idat_45;
  reg return_rsci_idat_44;
  reg return_rsci_idat_43;
  reg return_rsci_idat_42;
  reg return_rsci_idat_41;
  reg return_rsci_idat_40;
  reg return_rsci_idat_39;
  reg return_rsci_idat_38;
  reg return_rsci_idat_37;
  reg return_rsci_idat_36;
  reg return_rsci_idat_35;
  reg return_rsci_idat_34;
  reg return_rsci_idat_33;
  reg return_rsci_idat_32;
  reg return_rsci_idat_31;
  reg return_rsci_idat_30;
  reg return_rsci_idat_29;
  reg return_rsci_idat_28;
  reg return_rsci_idat_27;
  reg return_rsci_idat_26;
  reg return_rsci_idat_25;
  reg return_rsci_idat_24;
  reg return_rsci_idat_23;
  reg return_rsci_idat_22;
  reg return_rsci_idat_21;
  reg return_rsci_idat_20;
  reg return_rsci_idat_19;
  reg return_rsci_idat_18;
  reg return_rsci_idat_17;
  reg return_rsci_idat_16;
  reg return_rsci_idat_15;
  reg return_rsci_idat_14;
  reg return_rsci_idat_13;
  reg return_rsci_idat_12;
  reg return_rsci_idat_11;
  reg return_rsci_idat_10;
  reg return_rsci_idat_9;
  reg return_rsci_idat_8;
  reg return_rsci_idat_7;
  reg return_rsci_idat_6;
  reg return_rsci_idat_5;
  reg return_rsci_idat_4;
  reg return_rsci_idat_3;
  reg return_rsci_idat_2;
  reg return_rsci_idat_1;
  reg return_rsci_idat_0;
  wire [2:0] fsm_output;
  wire not_tmp_1;
  wire or_tmp_121;
  wire [4:0] i_3_4_0_sva_2;
  wire [5:0] nl_i_3_4_0_sva_2;
  reg [3:0] i_3_4_0_sva_3_0;
  reg reg_return_rsc_triosy_obj_ld_cse;
  reg L_15_sva;
  reg L_16_sva;
  reg L_14_sva;
  reg L_17_sva;
  reg L_13_sva;
  reg L_18_sva;
  reg L_12_sva;
  reg L_19_sva;
  reg L_11_sva;
  reg L_20_sva;
  reg L_10_sva;
  reg L_21_sva;
  reg L_9_sva;
  reg L_22_sva;
  reg L_8_sva;
  reg L_23_sva;
  reg L_7_sva;
  reg L_24_sva;
  reg L_6_sva;
  reg L_25_sva;
  reg L_5_sva;
  reg L_26_sva;
  reg L_4_sva;
  reg L_27_sva;
  reg L_3_sva;
  reg L_28_sva;
  reg L_2_sva;
  reg L_29_sva;
  reg L_1_sva;
  reg L_30_sva;
  reg L_0_sva;
  reg L_31_sva;
  reg R_15_sva;
  reg R_16_sva;
  reg R_14_sva;
  reg R_17_sva;
  reg R_13_sva;
  reg R_18_sva;
  reg R_12_sva;
  reg R_19_sva;
  reg R_11_sva;
  reg R_20_sva;
  reg R_10_sva;
  reg R_21_sva;
  reg R_9_sva;
  reg R_22_sva;
  reg R_8_sva;
  reg R_23_sva;
  reg R_7_sva;
  reg R_24_sva;
  reg R_6_sva;
  reg R_25_sva;
  reg R_5_sva;
  reg R_26_sva;
  reg R_4_sva;
  reg R_27_sva;
  reg R_3_sva;
  reg R_28_sva;
  reg R_2_sva;
  reg R_29_sva;
  reg R_1_sva;
  reg R_30_sva;
  reg R_0_sva;
  reg R_31_sva;
  reg C_1_13_sva;
  reg C_1_14_sva;
  reg C_1_12_sva;
  reg C_1_15_sva;
  reg C_1_11_sva;
  reg C_1_16_sva;
  reg C_1_10_sva;
  reg C_1_17_sva;
  reg C_1_9_sva;
  reg C_1_18_sva;
  reg C_1_8_sva;
  reg C_1_19_sva;
  reg C_1_7_sva;
  reg C_1_20_sva;
  reg C_1_6_sva;
  reg C_1_21_sva;
  reg C_1_5_sva;
  reg C_1_22_sva;
  reg C_1_4_sva;
  reg C_1_23_sva;
  reg C_1_3_sva;
  reg C_1_24_sva;
  reg C_1_2_sva;
  reg C_1_25_sva;
  reg C_1_1_sva;
  reg C_1_26_sva;
  reg C_1_0_sva;
  reg C_1_27_sva;
  reg D_1_13_sva;
  reg D_1_14_sva;
  reg D_1_12_sva;
  reg D_1_15_sva;
  reg D_1_11_sva;
  reg D_1_16_sva;
  reg D_1_10_sva;
  reg D_1_17_sva;
  reg D_1_9_sva;
  reg D_1_18_sva;
  reg D_1_8_sva;
  reg D_1_19_sva;
  reg D_1_7_sva;
  reg D_1_20_sva;
  reg D_1_6_sva;
  reg D_1_21_sva;
  reg D_1_5_sva;
  reg D_1_22_sva;
  reg D_1_4_sva;
  reg D_1_23_sva;
  reg D_1_3_sva;
  reg D_1_24_sva;
  reg D_1_2_sva;
  reg D_1_25_sva;
  reg D_1_1_sva;
  reg D_1_26_sva;
  reg D_1_0_sva;
  reg D_1_27_sva;
  wire R_24_sva_2;
  wire R_7_sva_2;
  wire R_16_sva_2;
  wire R_15_sva_2;
  wire R_8_sva_2;
  wire R_23_sva_2;
  wire R_0_sva_2;
  wire R_31_sva_2;
  wire R_25_sva_2;
  wire R_6_sva_2;
  wire R_17_sva_2;
  wire R_14_sva_2;
  wire R_9_sva_2;
  wire R_22_sva_2;
  wire R_1_sva_2;
  wire R_30_sva_2;
  wire R_26_sva_2;
  wire R_5_sva_2;
  wire R_18_sva_2;
  wire R_13_sva_2;
  wire R_10_sva_2;
  wire R_21_sva_2;
  wire R_2_sva_2;
  wire R_29_sva_2;
  wire R_27_sva_2;
  wire R_4_sva_2;
  wire R_19_sva_2;
  wire R_12_sva_2;
  wire R_11_sva_2;
  wire R_20_sva_2;
  wire R_3_sva_2;
  wire R_28_sva_2;
  wire D_1_26_sva_mx1;
  wire D_1_27_sva_mx1;
  wire D_1_0_sva_mx1;
  wire D_1_1_sva_mx1;
  wire D_1_3_sva_mx1;
  wire D_1_4_sva_mx1;
  wire D_1_5_sva_mx1;
  wire D_1_6_sva_mx1;
  wire D_1_7_sva_mx1;
  wire D_1_8_sva_mx1;
  wire D_1_9_sva_mx1;
  wire D_1_10_sva_mx1;
  wire D_1_11_sva_mx1;
  wire D_1_12_sva_mx1;
  wire D_1_14_sva_mx1;
  wire D_1_15_sva_mx1;
  wire D_1_16_sva_mx1;
  wire D_1_17_sva_mx1;
  wire D_1_19_sva_mx1;
  wire D_1_20_sva_mx1;
  wire D_1_22_sva_mx1;
  wire D_1_23_sva_mx1;
  wire D_1_24_sva_mx1;
  wire D_1_25_sva_mx1;
  wire C_1_26_sva_mx1;
  wire C_1_27_sva_mx1;
  wire C_1_0_sva_mx1;
  wire C_1_1_sva_mx1;
  wire C_1_2_sva_mx1;
  wire C_1_4_sva_mx1;
  wire C_1_5_sva_mx1;
  wire C_1_7_sva_mx1;
  wire C_1_8_sva_mx1;
  wire C_1_9_sva_mx1;
  wire C_1_11_sva_mx1;
  wire C_1_12_sva_mx1;
  wire C_1_13_sva_mx1;
  wire C_1_14_sva_mx1;
  wire C_1_15_sva_mx1;
  wire C_1_16_sva_mx1;
  wire C_1_17_sva_mx1;
  wire C_1_18_sva_mx1;
  wire C_1_20_sva_mx1;
  wire C_1_21_sva_mx1;
  wire C_1_22_sva_mx1;
  wire C_1_23_sva_mx1;
  wire C_1_24_sva_mx1;
  wire C_1_25_sva_mx1;
  wire [3:0] ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_1;
  wire [3:0] ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_1;
  wire [3:0] ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_1;
  wire [3:0] ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_1;
  wire [3:0] ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_1;
  wire [3:0] ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_1;
  wire [3:0] ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_1;
  wire [3:0] ROM_1i6_1o4_ce1b43b29576509b87f48de0e64c68b52f_1;

  wire[0:0] D_mux_9_nl;
  wire[0:0] D_mux_31_nl;
  wire[0:0] D_mux_41_nl;
  wire[0:0] D_mux_47_nl;
  wire[0:0] C_mux_11_nl;
  wire[0:0] C_mux_17_nl;
  wire[0:0] C_mux_25_nl;
  wire[0:0] C_mux_43_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [63:0] nl_return_rsci_idat;
  assign nl_return_rsci_idat = {return_rsci_idat_63 , return_rsci_idat_62 , return_rsci_idat_61
      , return_rsci_idat_60 , return_rsci_idat_59 , return_rsci_idat_58 , return_rsci_idat_57
      , return_rsci_idat_56 , return_rsci_idat_55 , return_rsci_idat_54 , return_rsci_idat_53
      , return_rsci_idat_52 , return_rsci_idat_51 , return_rsci_idat_50 , return_rsci_idat_49
      , return_rsci_idat_48 , return_rsci_idat_47 , return_rsci_idat_46 , return_rsci_idat_45
      , return_rsci_idat_44 , return_rsci_idat_43 , return_rsci_idat_42 , return_rsci_idat_41
      , return_rsci_idat_40 , return_rsci_idat_39 , return_rsci_idat_38 , return_rsci_idat_37
      , return_rsci_idat_36 , return_rsci_idat_35 , return_rsci_idat_34 , return_rsci_idat_33
      , return_rsci_idat_32 , return_rsci_idat_31 , return_rsci_idat_30 , return_rsci_idat_29
      , return_rsci_idat_28 , return_rsci_idat_27 , return_rsci_idat_26 , return_rsci_idat_25
      , return_rsci_idat_24 , return_rsci_idat_23 , return_rsci_idat_22 , return_rsci_idat_21
      , return_rsci_idat_20 , return_rsci_idat_19 , return_rsci_idat_18 , return_rsci_idat_17
      , return_rsci_idat_16 , return_rsci_idat_15 , return_rsci_idat_14 , return_rsci_idat_13
      , return_rsci_idat_12 , return_rsci_idat_11 , return_rsci_idat_10 , return_rsci_idat_9
      , return_rsci_idat_8 , return_rsci_idat_7 , return_rsci_idat_6 , return_rsci_idat_5
      , return_rsci_idat_4 , return_rsci_idat_3 , return_rsci_idat_2 , return_rsci_idat_1
      , return_rsci_idat_0};
  wire[0:0] loop_DES_rounds_xor_74_nl;
  wire[0:0] loop_DES_rounds_xor_79_nl;
  wire[0:0] loop_DES_rounds_xor_75_nl;
  wire[0:0] loop_DES_rounds_xor_76_nl;
  wire[0:0] loop_DES_rounds_xor_77_nl;
  wire[0:0] loop_DES_rounds_xor_78_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_rg_I_1;
  assign loop_DES_rounds_xor_74_nl = R_4_sva ^ D_1_10_sva_mx1;
  assign loop_DES_rounds_xor_79_nl = R_31_sva ^ D_1_24_sva_mx1;
  assign loop_DES_rounds_xor_75_nl = R_3_sva ^ D_1_14_sva_mx1;
  assign loop_DES_rounds_xor_76_nl = R_2_sva ^ D_1_6_sva_mx1;
  assign loop_DES_rounds_xor_77_nl = R_1_sva ^ D_1_20_sva_mx1;
  assign loop_DES_rounds_xor_78_nl = R_0_sva ^ D_1_27_sva_mx1;
  assign nl_U_ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_rg_I_1 = {loop_DES_rounds_xor_74_nl
      , loop_DES_rounds_xor_79_nl , loop_DES_rounds_xor_75_nl , loop_DES_rounds_xor_76_nl
      , loop_DES_rounds_xor_77_nl , loop_DES_rounds_xor_78_nl};
  wire[0:0] loop_DES_rounds_xor_50_nl;
  wire[0:0] loop_DES_rounds_xor_55_nl;
  wire[0:0] loop_DES_rounds_xor_51_nl;
  wire[0:0] loop_DES_rounds_xor_52_nl;
  wire[0:0] loop_DES_rounds_xor_53_nl;
  wire[0:0] loop_DES_rounds_xor_54_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_rg_I_1;
  assign loop_DES_rounds_xor_50_nl = R_20_sva ^ C_1_12_sva_mx1;
  assign loop_DES_rounds_xor_55_nl = R_15_sva ^ C_1_26_sva_mx1;
  assign loop_DES_rounds_xor_51_nl = R_19_sva ^ C_1_21_sva_mx1;
  assign loop_DES_rounds_xor_52_nl = R_18_sva ^ C_1_1_sva_mx1;
  assign loop_DES_rounds_xor_53_nl = R_17_sva ^ C_1_8_sva_mx1;
  assign loop_DES_rounds_xor_54_nl = R_16_sva ^ C_1_15_sva_mx1;
  assign nl_U_ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_rg_I_1 = {loop_DES_rounds_xor_50_nl
      , loop_DES_rounds_xor_55_nl , loop_DES_rounds_xor_51_nl , loop_DES_rounds_xor_52_nl
      , loop_DES_rounds_xor_53_nl , loop_DES_rounds_xor_54_nl};
  wire[0:0] loop_DES_rounds_xor_68_nl;
  wire[0:0] loop_DES_rounds_xor_73_nl;
  wire[0:0] loop_DES_rounds_xor_69_nl;
  wire[0:0] loop_DES_rounds_xor_70_nl;
  wire[0:0] loop_DES_rounds_xor_71_nl;
  wire[0:0] loop_DES_rounds_xor_72_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_rg_I_1;
  assign loop_DES_rounds_xor_68_nl = R_8_sva ^ D_1_12_sva_mx1;
  assign loop_DES_rounds_xor_73_nl = R_3_sva ^ D_1_3_sva_mx1;
  assign loop_DES_rounds_xor_69_nl = R_7_sva ^ D_1_7_sva_mx1;
  assign loop_DES_rounds_xor_70_nl = R_6_sva ^ D_1_17_sva_mx1;
  assign loop_DES_rounds_xor_71_nl = R_5_sva ^ D_1_0_sva_mx1;
  assign loop_DES_rounds_xor_72_nl = R_4_sva ^ D_1_22_sva_mx1;
  assign nl_U_ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_rg_I_1 = {loop_DES_rounds_xor_68_nl
      , loop_DES_rounds_xor_73_nl , loop_DES_rounds_xor_69_nl , loop_DES_rounds_xor_70_nl
      , loop_DES_rounds_xor_71_nl , loop_DES_rounds_xor_72_nl};
  wire[0:0] loop_DES_rounds_xor_44_nl;
  wire[0:0] loop_DES_rounds_xor_49_nl;
  wire[0:0] loop_DES_rounds_xor_45_nl;
  wire[0:0] loop_DES_rounds_xor_46_nl;
  wire[0:0] loop_DES_rounds_xor_47_nl;
  wire[0:0] loop_DES_rounds_xor_48_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_rg_I_1;
  assign loop_DES_rounds_xor_44_nl = R_24_sva ^ C_1_5_sva_mx1;
  assign loop_DES_rounds_xor_49_nl = R_19_sva ^ C_1_20_sva_mx1;
  assign loop_DES_rounds_xor_45_nl = R_23_sva ^ C_1_9_sva_mx1;
  assign loop_DES_rounds_xor_46_nl = R_22_sva ^ C_1_16_sva_mx1;
  assign loop_DES_rounds_xor_47_nl = R_21_sva ^ C_1_24_sva_mx1;
  assign loop_DES_rounds_xor_48_nl = R_20_sva ^ C_1_2_sva_mx1;
  assign nl_U_ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_rg_I_1 = {loop_DES_rounds_xor_44_nl
      , loop_DES_rounds_xor_49_nl , loop_DES_rounds_xor_45_nl , loop_DES_rounds_xor_46_nl
      , loop_DES_rounds_xor_47_nl , loop_DES_rounds_xor_48_nl};
  wire[0:0] loop_DES_rounds_xor_62_nl;
  wire[0:0] loop_DES_rounds_xor_67_nl;
  wire[0:0] loop_DES_rounds_xor_63_nl;
  wire[0:0] loop_DES_rounds_xor_64_nl;
  wire[0:0] loop_DES_rounds_xor_65_nl;
  wire[0:0] loop_DES_rounds_xor_66_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_rg_I_1;
  assign loop_DES_rounds_xor_62_nl = R_12_sva ^ D_1_26_sva_mx1;
  assign loop_DES_rounds_xor_67_nl = R_7_sva ^ D_1_8_sva_mx1;
  assign loop_DES_rounds_xor_63_nl = R_11_sva ^ D_1_16_sva_mx1;
  assign loop_DES_rounds_xor_64_nl = R_10_sva ^ D_1_5_sva_mx1;
  assign loop_DES_rounds_xor_65_nl = R_9_sva ^ D_1_11_sva_mx1;
  assign loop_DES_rounds_xor_66_nl = R_8_sva ^ D_1_23_sva_mx1;
  assign nl_U_ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_rg_I_1 = {loop_DES_rounds_xor_62_nl
      , loop_DES_rounds_xor_67_nl , loop_DES_rounds_xor_63_nl , loop_DES_rounds_xor_64_nl
      , loop_DES_rounds_xor_65_nl , loop_DES_rounds_xor_66_nl};
  wire[0:0] loop_DES_rounds_xor_38_nl;
  wire[0:0] loop_DES_rounds_xor_43_nl;
  wire[0:0] loop_DES_rounds_xor_39_nl;
  wire[0:0] loop_DES_rounds_xor_40_nl;
  wire[0:0] loop_DES_rounds_xor_41_nl;
  wire[0:0] loop_DES_rounds_xor_42_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_rg_I_1;
  assign loop_DES_rounds_xor_38_nl = R_28_sva ^ C_1_25_sva_mx1;
  assign loop_DES_rounds_xor_43_nl = R_23_sva ^ C_1_18_sva_mx1;
  assign loop_DES_rounds_xor_39_nl = R_27_sva ^ C_1_0_sva_mx1;
  assign loop_DES_rounds_xor_40_nl = R_26_sva ^ C_1_13_sva_mx1;
  assign loop_DES_rounds_xor_41_nl = R_25_sva ^ C_1_22_sva_mx1;
  assign loop_DES_rounds_xor_42_nl = R_24_sva ^ C_1_7_sva_mx1;
  assign nl_U_ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_rg_I_1 = {loop_DES_rounds_xor_38_nl
      , loop_DES_rounds_xor_43_nl , loop_DES_rounds_xor_39_nl , loop_DES_rounds_xor_40_nl
      , loop_DES_rounds_xor_41_nl , loop_DES_rounds_xor_42_nl};
  wire[0:0] loop_DES_rounds_xor_56_nl;
  wire[0:0] loop_DES_rounds_xor_61_nl;
  wire[0:0] loop_DES_rounds_xor_57_nl;
  wire[0:0] loop_DES_rounds_xor_58_nl;
  wire[0:0] loop_DES_rounds_xor_59_nl;
  wire[0:0] loop_DES_rounds_xor_60_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_rg_I_1;
  assign loop_DES_rounds_xor_56_nl = R_16_sva ^ D_1_15_sva_mx1;
  assign loop_DES_rounds_xor_61_nl = R_11_sva ^ D_1_1_sva_mx1;
  assign loop_DES_rounds_xor_57_nl = R_15_sva ^ D_1_4_sva_mx1;
  assign loop_DES_rounds_xor_58_nl = R_14_sva ^ D_1_25_sva_mx1;
  assign loop_DES_rounds_xor_59_nl = R_13_sva ^ D_1_19_sva_mx1;
  assign loop_DES_rounds_xor_60_nl = R_12_sva ^ D_1_9_sva_mx1;
  assign nl_U_ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_rg_I_1 = {loop_DES_rounds_xor_56_nl
      , loop_DES_rounds_xor_61_nl , loop_DES_rounds_xor_57_nl , loop_DES_rounds_xor_58_nl
      , loop_DES_rounds_xor_59_nl , loop_DES_rounds_xor_60_nl};
  wire[0:0] loop_DES_rounds_xor_nl;
  wire[0:0] loop_DES_rounds_xor_37_nl;
  wire[0:0] loop_DES_rounds_xor_33_nl;
  wire[0:0] loop_DES_rounds_xor_34_nl;
  wire[0:0] loop_DES_rounds_xor_35_nl;
  wire[0:0] loop_DES_rounds_xor_36_nl;
  wire [5:0] nl_U_ROM_1i6_1o4_ce1b43b29576509b87f48de0e64c68b52f_rg_I_1;
  assign loop_DES_rounds_xor_nl = R_0_sva ^ C_1_14_sva_mx1;
  assign loop_DES_rounds_xor_37_nl = R_27_sva ^ C_1_23_sva_mx1;
  assign loop_DES_rounds_xor_33_nl = R_31_sva ^ C_1_11_sva_mx1;
  assign loop_DES_rounds_xor_34_nl = R_30_sva ^ C_1_17_sva_mx1;
  assign loop_DES_rounds_xor_35_nl = R_29_sva ^ C_1_4_sva_mx1;
  assign loop_DES_rounds_xor_36_nl = R_28_sva ^ C_1_27_sva_mx1;
  assign nl_U_ROM_1i6_1o4_ce1b43b29576509b87f48de0e64c68b52f_rg_I_1 = {loop_DES_rounds_xor_nl
      , loop_DES_rounds_xor_37_nl , loop_DES_rounds_xor_33_nl , loop_DES_rounds_xor_34_nl
      , loop_DES_rounds_xor_35_nl , loop_DES_rounds_xor_36_nl};
  wire [0:0] nl_des_check_core_core_fsm_inst_loop_DES_rounds_C_0_tr0;
  assign nl_des_check_core_core_fsm_inst_loop_DES_rounds_C_0_tr0 = i_3_4_0_sva_2[4];
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd64)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd64)) key_rsci (
      .dat(key_rsc_dat),
      .idat(key_rsci_idat)
    );
  ccs_out_v1 #(.rscid(32'sd3),
  .width(32'sd64)) return_rsci (
      .idat(nl_return_rsci_idat[63:0]),
      .dat(return_rsc_dat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) input_rsc_triosy_obj (
      .ld(reg_return_rsc_triosy_obj_ld_cse),
      .lz(input_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) key_rsc_triosy_obj (
      .ld(reg_return_rsc_triosy_obj_ld_cse),
      .lz(key_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) return_rsc_triosy_obj (
      .ld(reg_return_rsc_triosy_obj_ld_cse),
      .lz(return_rsc_triosy_lz)
    );
  ROM_1i6_1o4_ef4da7ff735c86ba85f23e51741d972cb3  U_ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_1)
    );
  ROM_1i6_1o4_d0e242163cbb0b2ce9c4399bc1cb50f5b3  U_ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_1)
    );
  ROM_1i6_1o4_752c7ca65a598ada4acee0cd63d199c3b3  U_ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_1)
    );
  ROM_1i6_1o4_3c5c29b75c561d2b741f22e5a3a569dbb3  U_ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_1)
    );
  ROM_1i6_1o4_51ba7157b272cd3b87451219caf38e7cb3  U_ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_1)
    );
  ROM_1i6_1o4_cfafff97e973ca9580e646fecdc2f814b3  U_ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_1)
    );
  ROM_1i6_1o4_ef717c7c87dc90ac6f7b34d533fe115fb3  U_ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_1)
    );
  ROM_1i6_1o4_8f60b2fc4a3ee4cef30040071bc0219cb3  U_ROM_1i6_1o4_ce1b43b29576509b87f48de0e64c68b52f_rg
      (
      .I_1(nl_U_ROM_1i6_1o4_ce1b43b29576509b87f48de0e64c68b52f_rg_I_1[5:0]),
      .O_1(ROM_1i6_1o4_ce1b43b29576509b87f48de0e64c68b52f_1)
    );
  des_check_core_core_fsm des_check_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .loop_DES_rounds_C_0_tr0(nl_des_check_core_core_fsm_inst_loop_DES_rounds_C_0_tr0[0:0])
    );
  assign R_24_sva_2 = L_24_sva ^ (ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_1[3]);
  assign R_7_sva_2 = L_7_sva ^ (ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_1[1]);
  assign R_16_sva_2 = L_16_sva ^ (ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_1[2]);
  assign R_15_sva_2 = L_15_sva ^ (ROM_1i6_1o4_ce1b43b29576509b87f48de0e64c68b52f_1[2]);
  assign R_8_sva_2 = L_8_sva ^ (ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_1[3]);
  assign R_23_sva_2 = L_23_sva ^ (ROM_1i6_1o4_ce1b43b29576509b87f48de0e64c68b52f_1[3]);
  assign R_0_sva_2 = L_0_sva ^ (ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_1[3]);
  assign R_31_sva_2 = L_31_sva ^ (ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_1[0]);
  assign R_25_sva_2 = L_25_sva ^ (ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_1[0]);
  assign R_6_sva_2 = L_6_sva ^ (ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_1[3]);
  assign R_17_sva_2 = L_17_sva ^ (ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_1[1]);
  assign R_14_sva_2 = L_14_sva ^ (ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_1[0]);
  assign R_9_sva_2 = L_9_sva ^ (ROM_1i6_1o4_ce1b43b29576509b87f48de0e64c68b52f_1[1]);
  assign R_22_sva_2 = L_22_sva ^ (ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_1[1]);
  assign R_1_sva_2 = L_1_sva ^ (ROM_1i6_1o4_ce1b43b29576509b87f48de0e64c68b52f_1[0]);
  assign R_30_sva_2 = L_30_sva ^ (ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_1[1]);
  assign R_26_sva_2 = L_26_sva ^ (ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_1[0]);
  assign R_5_sva_2 = L_5_sva ^ (ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_1[2]);
  assign R_18_sva_2 = L_18_sva ^ (ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_1[2]);
  assign R_13_sva_2 = L_13_sva ^ (ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_1[0]);
  assign R_10_sva_2 = L_10_sva ^ (ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_1[1]);
  assign R_21_sva_2 = L_21_sva ^ (ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_1[1]);
  assign R_2_sva_2 = L_2_sva ^ (ROM_1i6_1o4_644850663d96c9b3c8a27f69784ee5782f_1[1]);
  assign R_29_sva_2 = L_29_sva ^ (ROM_1i6_1o4_5d76c79e05be4dd136865bde1aaf01c82f_1[0]);
  assign R_27_sva_2 = L_27_sva ^ (ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_1[3]);
  assign R_4_sva_2 = L_4_sva ^ (ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_1[2]);
  assign R_19_sva_2 = L_19_sva ^ (ROM_1i6_1o4_79fefe0558b80605fe451e50421a35632f_1[3]);
  assign R_12_sva_2 = L_12_sva ^ (ROM_1i6_1o4_573cd39ad7d789c17a1aa9155f1a1a9b2f_1[2]);
  assign R_11_sva_2 = L_11_sva ^ (ROM_1i6_1o4_35be3ef31c93661f5e99f6752adf3f622f_1[0]);
  assign R_20_sva_2 = L_20_sva ^ (ROM_1i6_1o4_dcd0439231154fad8f91fc0951bedbc32f_1[2]);
  assign R_3_sva_2 = L_3_sva ^ (ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_1[2]);
  assign R_28_sva_2 = L_28_sva ^ (ROM_1i6_1o4_67cbe7fa3f0828c413079bd7c0dc864f2f_1[3]);
  assign D_1_26_sva_mx1 = MUX_s_1_2_2(D_1_25_sva, D_1_24_sva, not_tmp_1);
  assign D_1_27_sva_mx1 = MUX_s_1_2_2(D_1_26_sva, D_1_25_sva, not_tmp_1);
  assign D_1_0_sva_mx1 = MUX_s_1_2_2(D_1_27_sva, D_1_26_sva, not_tmp_1);
  assign D_1_1_sva_mx1 = MUX_s_1_2_2(D_1_0_sva, D_1_27_sva, not_tmp_1);
  assign D_1_3_sva_mx1 = MUX_s_1_2_2(D_1_2_sva, D_1_1_sva, not_tmp_1);
  assign D_1_4_sva_mx1 = MUX_s_1_2_2(D_1_3_sva, D_1_2_sva, not_tmp_1);
  assign D_1_5_sva_mx1 = MUX_s_1_2_2(D_1_4_sva, D_1_3_sva, not_tmp_1);
  assign D_1_6_sva_mx1 = MUX_s_1_2_2(D_1_5_sva, D_1_4_sva, not_tmp_1);
  assign D_1_7_sva_mx1 = MUX_s_1_2_2(D_1_6_sva, D_1_5_sva, not_tmp_1);
  assign D_1_8_sva_mx1 = MUX_s_1_2_2(D_1_7_sva, D_1_6_sva, not_tmp_1);
  assign D_1_9_sva_mx1 = MUX_s_1_2_2(D_1_8_sva, D_1_7_sva, not_tmp_1);
  assign D_1_10_sva_mx1 = MUX_s_1_2_2(D_1_9_sva, D_1_8_sva, not_tmp_1);
  assign D_1_11_sva_mx1 = MUX_s_1_2_2(D_1_10_sva, D_1_9_sva, not_tmp_1);
  assign D_1_12_sva_mx1 = MUX_s_1_2_2(D_1_11_sva, D_1_10_sva, not_tmp_1);
  assign D_1_14_sva_mx1 = MUX_s_1_2_2(D_1_13_sva, D_1_12_sva, not_tmp_1);
  assign D_1_15_sva_mx1 = MUX_s_1_2_2(D_1_14_sva, D_1_13_sva, not_tmp_1);
  assign D_1_16_sva_mx1 = MUX_s_1_2_2(D_1_15_sva, D_1_14_sva, not_tmp_1);
  assign D_1_17_sva_mx1 = MUX_s_1_2_2(D_1_16_sva, D_1_15_sva, not_tmp_1);
  assign D_1_19_sva_mx1 = MUX_s_1_2_2(D_1_18_sva, D_1_17_sva, not_tmp_1);
  assign D_1_20_sva_mx1 = MUX_s_1_2_2(D_1_19_sva, D_1_18_sva, not_tmp_1);
  assign D_1_22_sva_mx1 = MUX_s_1_2_2(D_1_21_sva, D_1_20_sva, not_tmp_1);
  assign D_1_23_sva_mx1 = MUX_s_1_2_2(D_1_22_sva, D_1_21_sva, not_tmp_1);
  assign D_1_24_sva_mx1 = MUX_s_1_2_2(D_1_23_sva, D_1_22_sva, not_tmp_1);
  assign D_1_25_sva_mx1 = MUX_s_1_2_2(D_1_24_sva, D_1_23_sva, not_tmp_1);
  assign C_1_26_sva_mx1 = MUX_s_1_2_2(C_1_25_sva, C_1_24_sva, not_tmp_1);
  assign C_1_27_sva_mx1 = MUX_s_1_2_2(C_1_26_sva, C_1_25_sva, not_tmp_1);
  assign C_1_0_sva_mx1 = MUX_s_1_2_2(C_1_27_sva, C_1_26_sva, not_tmp_1);
  assign C_1_1_sva_mx1 = MUX_s_1_2_2(C_1_0_sva, C_1_27_sva, not_tmp_1);
  assign C_1_2_sva_mx1 = MUX_s_1_2_2(C_1_1_sva, C_1_0_sva, not_tmp_1);
  assign C_1_4_sva_mx1 = MUX_s_1_2_2(C_1_3_sva, C_1_2_sva, not_tmp_1);
  assign C_1_5_sva_mx1 = MUX_s_1_2_2(C_1_4_sva, C_1_3_sva, not_tmp_1);
  assign C_1_7_sva_mx1 = MUX_s_1_2_2(C_1_6_sva, C_1_5_sva, not_tmp_1);
  assign C_1_8_sva_mx1 = MUX_s_1_2_2(C_1_7_sva, C_1_6_sva, not_tmp_1);
  assign C_1_9_sva_mx1 = MUX_s_1_2_2(C_1_8_sva, C_1_7_sva, not_tmp_1);
  assign C_1_11_sva_mx1 = MUX_s_1_2_2(C_1_10_sva, C_1_9_sva, not_tmp_1);
  assign C_1_12_sva_mx1 = MUX_s_1_2_2(C_1_11_sva, C_1_10_sva, not_tmp_1);
  assign C_1_13_sva_mx1 = MUX_s_1_2_2(C_1_12_sva, C_1_11_sva, not_tmp_1);
  assign C_1_14_sva_mx1 = MUX_s_1_2_2(C_1_13_sva, C_1_12_sva, not_tmp_1);
  assign C_1_15_sva_mx1 = MUX_s_1_2_2(C_1_14_sva, C_1_13_sva, not_tmp_1);
  assign C_1_16_sva_mx1 = MUX_s_1_2_2(C_1_15_sva, C_1_14_sva, not_tmp_1);
  assign C_1_17_sva_mx1 = MUX_s_1_2_2(C_1_16_sva, C_1_15_sva, not_tmp_1);
  assign C_1_18_sva_mx1 = MUX_s_1_2_2(C_1_17_sva, C_1_16_sva, not_tmp_1);
  assign C_1_20_sva_mx1 = MUX_s_1_2_2(C_1_19_sva, C_1_18_sva, not_tmp_1);
  assign C_1_21_sva_mx1 = MUX_s_1_2_2(C_1_20_sva, C_1_19_sva, not_tmp_1);
  assign C_1_22_sva_mx1 = MUX_s_1_2_2(C_1_21_sva, C_1_20_sva, not_tmp_1);
  assign C_1_23_sva_mx1 = MUX_s_1_2_2(C_1_22_sva, C_1_21_sva, not_tmp_1);
  assign C_1_24_sva_mx1 = MUX_s_1_2_2(C_1_23_sva, C_1_22_sva, not_tmp_1);
  assign C_1_25_sva_mx1 = MUX_s_1_2_2(C_1_24_sva, C_1_23_sva, not_tmp_1);
  assign nl_i_3_4_0_sva_2 = conv_u2s_4_5(i_3_4_0_sva_3_0) + 5'b00001;
  assign i_3_4_0_sva_2 = nl_i_3_4_0_sva_2[4:0];
  assign not_tmp_1 = ~(((i_3_4_0_sva_3_0==4'b1111)) | ((i_3_4_0_sva_3_0==4'b1000))
      | (~((~((i_3_4_0_sva_3_0==4'b0001))) & ((i_3_4_0_sva_3_0!=4'b0000)))));
  assign or_tmp_121 = ~((i_3_4_0_sva_2[4]) & (fsm_output[1]));
  always @(posedge clk) begin
    if ( rst ) begin
      R_24_sva <= 1'b0;
      R_7_sva <= 1'b0;
      R_16_sva <= 1'b0;
      R_15_sva <= 1'b0;
      R_8_sva <= 1'b0;
      R_23_sva <= 1'b0;
      R_0_sva <= 1'b0;
      R_31_sva <= 1'b0;
      R_25_sva <= 1'b0;
      R_6_sva <= 1'b0;
      R_17_sva <= 1'b0;
      R_14_sva <= 1'b0;
      R_9_sva <= 1'b0;
      R_22_sva <= 1'b0;
      R_1_sva <= 1'b0;
      R_30_sva <= 1'b0;
      R_26_sva <= 1'b0;
      R_5_sva <= 1'b0;
      R_18_sva <= 1'b0;
      R_13_sva <= 1'b0;
      R_10_sva <= 1'b0;
      R_21_sva <= 1'b0;
      R_2_sva <= 1'b0;
      R_29_sva <= 1'b0;
      R_27_sva <= 1'b0;
      R_4_sva <= 1'b0;
      R_19_sva <= 1'b0;
      R_12_sva <= 1'b0;
      R_11_sva <= 1'b0;
      R_20_sva <= 1'b0;
      R_3_sva <= 1'b0;
      R_28_sva <= 1'b0;
      i_3_4_0_sva_3_0 <= 4'b0000;
      L_31_sva <= 1'b0;
      L_0_sva <= 1'b0;
      L_30_sva <= 1'b0;
      L_1_sva <= 1'b0;
      L_29_sva <= 1'b0;
      L_2_sva <= 1'b0;
      L_28_sva <= 1'b0;
      L_3_sva <= 1'b0;
      L_27_sva <= 1'b0;
      L_4_sva <= 1'b0;
      L_26_sva <= 1'b0;
      L_5_sva <= 1'b0;
      L_25_sva <= 1'b0;
      L_6_sva <= 1'b0;
      L_24_sva <= 1'b0;
      L_7_sva <= 1'b0;
      L_23_sva <= 1'b0;
      L_8_sva <= 1'b0;
      L_22_sva <= 1'b0;
      L_9_sva <= 1'b0;
      L_21_sva <= 1'b0;
      L_10_sva <= 1'b0;
      L_20_sva <= 1'b0;
      L_11_sva <= 1'b0;
      L_19_sva <= 1'b0;
      L_12_sva <= 1'b0;
      L_18_sva <= 1'b0;
      L_13_sva <= 1'b0;
      L_17_sva <= 1'b0;
      L_14_sva <= 1'b0;
      L_16_sva <= 1'b0;
      L_15_sva <= 1'b0;
      D_1_26_sva <= 1'b0;
      D_1_27_sva <= 1'b0;
      D_1_0_sva <= 1'b0;
      D_1_1_sva <= 1'b0;
      D_1_2_sva <= 1'b0;
      D_1_3_sva <= 1'b0;
      D_1_4_sva <= 1'b0;
      D_1_5_sva <= 1'b0;
      D_1_6_sva <= 1'b0;
      D_1_7_sva <= 1'b0;
      D_1_8_sva <= 1'b0;
      D_1_9_sva <= 1'b0;
      D_1_10_sva <= 1'b0;
      D_1_11_sva <= 1'b0;
      D_1_12_sva <= 1'b0;
      D_1_13_sva <= 1'b0;
      D_1_14_sva <= 1'b0;
      D_1_15_sva <= 1'b0;
      D_1_16_sva <= 1'b0;
      D_1_17_sva <= 1'b0;
      D_1_18_sva <= 1'b0;
      D_1_19_sva <= 1'b0;
      D_1_20_sva <= 1'b0;
      D_1_21_sva <= 1'b0;
      D_1_22_sva <= 1'b0;
      D_1_23_sva <= 1'b0;
      D_1_24_sva <= 1'b0;
      D_1_25_sva <= 1'b0;
      C_1_26_sva <= 1'b0;
      C_1_27_sva <= 1'b0;
      C_1_0_sva <= 1'b0;
      C_1_1_sva <= 1'b0;
      C_1_2_sva <= 1'b0;
      C_1_3_sva <= 1'b0;
      C_1_4_sva <= 1'b0;
      C_1_5_sva <= 1'b0;
      C_1_6_sva <= 1'b0;
      C_1_7_sva <= 1'b0;
      C_1_8_sva <= 1'b0;
      C_1_9_sva <= 1'b0;
      C_1_10_sva <= 1'b0;
      C_1_11_sva <= 1'b0;
      C_1_12_sva <= 1'b0;
      C_1_13_sva <= 1'b0;
      C_1_14_sva <= 1'b0;
      C_1_15_sva <= 1'b0;
      C_1_16_sva <= 1'b0;
      C_1_17_sva <= 1'b0;
      C_1_18_sva <= 1'b0;
      C_1_19_sva <= 1'b0;
      C_1_20_sva <= 1'b0;
      C_1_21_sva <= 1'b0;
      C_1_22_sva <= 1'b0;
      C_1_23_sva <= 1'b0;
      C_1_24_sva <= 1'b0;
      C_1_25_sva <= 1'b0;
      reg_return_rsc_triosy_obj_ld_cse <= 1'b0;
    end
    else begin
      R_24_sva <= MUX_s_1_2_2((input_rsci_idat[63]), R_24_sva_2, fsm_output[1]);
      R_7_sva <= MUX_s_1_2_2((input_rsci_idat[1]), R_7_sva_2, fsm_output[1]);
      R_16_sva <= MUX_s_1_2_2((input_rsci_idat[61]), R_16_sva_2, fsm_output[1]);
      R_15_sva <= MUX_s_1_2_2((input_rsci_idat[3]), R_15_sva_2, fsm_output[1]);
      R_8_sva <= MUX_s_1_2_2((input_rsci_idat[59]), R_8_sva_2, fsm_output[1]);
      R_23_sva <= MUX_s_1_2_2((input_rsci_idat[5]), R_23_sva_2, fsm_output[1]);
      R_0_sva <= MUX_s_1_2_2((input_rsci_idat[57]), R_0_sva_2, fsm_output[1]);
      R_31_sva <= MUX_s_1_2_2((input_rsci_idat[7]), R_31_sva_2, fsm_output[1]);
      R_25_sva <= MUX_s_1_2_2((input_rsci_idat[55]), R_25_sva_2, fsm_output[1]);
      R_6_sva <= MUX_s_1_2_2((input_rsci_idat[9]), R_6_sva_2, fsm_output[1]);
      R_17_sva <= MUX_s_1_2_2((input_rsci_idat[53]), R_17_sva_2, fsm_output[1]);
      R_14_sva <= MUX_s_1_2_2((input_rsci_idat[11]), R_14_sva_2, fsm_output[1]);
      R_9_sva <= MUX_s_1_2_2((input_rsci_idat[51]), R_9_sva_2, fsm_output[1]);
      R_22_sva <= MUX_s_1_2_2((input_rsci_idat[13]), R_22_sva_2, fsm_output[1]);
      R_1_sva <= MUX_s_1_2_2((input_rsci_idat[49]), R_1_sva_2, fsm_output[1]);
      R_30_sva <= MUX_s_1_2_2((input_rsci_idat[15]), R_30_sva_2, fsm_output[1]);
      R_26_sva <= MUX_s_1_2_2((input_rsci_idat[47]), R_26_sva_2, fsm_output[1]);
      R_5_sva <= MUX_s_1_2_2((input_rsci_idat[17]), R_5_sva_2, fsm_output[1]);
      R_18_sva <= MUX_s_1_2_2((input_rsci_idat[45]), R_18_sva_2, fsm_output[1]);
      R_13_sva <= MUX_s_1_2_2((input_rsci_idat[19]), R_13_sva_2, fsm_output[1]);
      R_10_sva <= MUX_s_1_2_2((input_rsci_idat[43]), R_10_sva_2, fsm_output[1]);
      R_21_sva <= MUX_s_1_2_2((input_rsci_idat[21]), R_21_sva_2, fsm_output[1]);
      R_2_sva <= MUX_s_1_2_2((input_rsci_idat[41]), R_2_sva_2, fsm_output[1]);
      R_29_sva <= MUX_s_1_2_2((input_rsci_idat[23]), R_29_sva_2, fsm_output[1]);
      R_27_sva <= MUX_s_1_2_2((input_rsci_idat[39]), R_27_sva_2, fsm_output[1]);
      R_4_sva <= MUX_s_1_2_2((input_rsci_idat[25]), R_4_sva_2, fsm_output[1]);
      R_19_sva <= MUX_s_1_2_2((input_rsci_idat[37]), R_19_sva_2, fsm_output[1]);
      R_12_sva <= MUX_s_1_2_2((input_rsci_idat[27]), R_12_sva_2, fsm_output[1]);
      R_11_sva <= MUX_s_1_2_2((input_rsci_idat[35]), R_11_sva_2, fsm_output[1]);
      R_20_sva <= MUX_s_1_2_2((input_rsci_idat[29]), R_20_sva_2, fsm_output[1]);
      R_3_sva <= MUX_s_1_2_2((input_rsci_idat[33]), R_3_sva_2, fsm_output[1]);
      R_28_sva <= MUX_s_1_2_2((input_rsci_idat[31]), R_28_sva_2, fsm_output[1]);
      i_3_4_0_sva_3_0 <= MUX_v_4_2_2(4'b0000, (i_3_4_0_sva_2[3:0]), (fsm_output[1]));
      L_31_sva <= MUX_s_1_2_2((input_rsci_idat[6]), R_31_sva, fsm_output[1]);
      L_0_sva <= MUX_s_1_2_2((input_rsci_idat[56]), R_0_sva, fsm_output[1]);
      L_30_sva <= MUX_s_1_2_2((input_rsci_idat[14]), R_30_sva, fsm_output[1]);
      L_1_sva <= MUX_s_1_2_2((input_rsci_idat[48]), R_1_sva, fsm_output[1]);
      L_29_sva <= MUX_s_1_2_2((input_rsci_idat[22]), R_29_sva, fsm_output[1]);
      L_2_sva <= MUX_s_1_2_2((input_rsci_idat[40]), R_2_sva, fsm_output[1]);
      L_28_sva <= MUX_s_1_2_2((input_rsci_idat[30]), R_28_sva, fsm_output[1]);
      L_3_sva <= MUX_s_1_2_2((input_rsci_idat[32]), R_3_sva, fsm_output[1]);
      L_27_sva <= MUX_s_1_2_2((input_rsci_idat[38]), R_27_sva, fsm_output[1]);
      L_4_sva <= MUX_s_1_2_2((input_rsci_idat[24]), R_4_sva, fsm_output[1]);
      L_26_sva <= MUX_s_1_2_2((input_rsci_idat[46]), R_26_sva, fsm_output[1]);
      L_5_sva <= MUX_s_1_2_2((input_rsci_idat[16]), R_5_sva, fsm_output[1]);
      L_25_sva <= MUX_s_1_2_2((input_rsci_idat[54]), R_25_sva, fsm_output[1]);
      L_6_sva <= MUX_s_1_2_2((input_rsci_idat[8]), R_6_sva, fsm_output[1]);
      L_24_sva <= MUX_s_1_2_2((input_rsci_idat[62]), R_24_sva, fsm_output[1]);
      L_7_sva <= MUX_s_1_2_2((input_rsci_idat[0]), R_7_sva, fsm_output[1]);
      L_23_sva <= MUX_s_1_2_2((input_rsci_idat[4]), R_23_sva, fsm_output[1]);
      L_8_sva <= MUX_s_1_2_2((input_rsci_idat[58]), R_8_sva, fsm_output[1]);
      L_22_sva <= MUX_s_1_2_2((input_rsci_idat[12]), R_22_sva, fsm_output[1]);
      L_9_sva <= MUX_s_1_2_2((input_rsci_idat[50]), R_9_sva, fsm_output[1]);
      L_21_sva <= MUX_s_1_2_2((input_rsci_idat[20]), R_21_sva, fsm_output[1]);
      L_10_sva <= MUX_s_1_2_2((input_rsci_idat[42]), R_10_sva, fsm_output[1]);
      L_20_sva <= MUX_s_1_2_2((input_rsci_idat[28]), R_20_sva, fsm_output[1]);
      L_11_sva <= MUX_s_1_2_2((input_rsci_idat[34]), R_11_sva, fsm_output[1]);
      L_19_sva <= MUX_s_1_2_2((input_rsci_idat[36]), R_19_sva, fsm_output[1]);
      L_12_sva <= MUX_s_1_2_2((input_rsci_idat[26]), R_12_sva, fsm_output[1]);
      L_18_sva <= MUX_s_1_2_2((input_rsci_idat[44]), R_18_sva, fsm_output[1]);
      L_13_sva <= MUX_s_1_2_2((input_rsci_idat[18]), R_13_sva, fsm_output[1]);
      L_17_sva <= MUX_s_1_2_2((input_rsci_idat[52]), R_17_sva, fsm_output[1]);
      L_14_sva <= MUX_s_1_2_2((input_rsci_idat[10]), R_14_sva, fsm_output[1]);
      L_16_sva <= MUX_s_1_2_2((input_rsci_idat[60]), R_16_sva, fsm_output[1]);
      L_15_sva <= MUX_s_1_2_2((input_rsci_idat[2]), R_15_sva, fsm_output[1]);
      D_1_26_sva <= MUX_s_1_2_2((key_rsci_idat[9]), D_1_26_sva_mx1, fsm_output[1]);
      D_1_27_sva <= MUX_s_1_2_2((key_rsci_idat[1]), D_1_27_sva_mx1, fsm_output[1]);
      D_1_0_sva <= MUX_s_1_2_2((key_rsci_idat[60]), D_1_0_sva_mx1, fsm_output[1]);
      D_1_1_sva <= MUX_s_1_2_2((key_rsci_idat[52]), D_1_1_sva_mx1, fsm_output[1]);
      D_1_2_sva <= MUX_s_1_2_2((key_rsci_idat[44]), D_mux_9_nl, fsm_output[1]);
      D_1_3_sva <= MUX_s_1_2_2((key_rsci_idat[36]), D_1_3_sva_mx1, fsm_output[1]);
      D_1_4_sva <= MUX_s_1_2_2((key_rsci_idat[59]), D_1_4_sva_mx1, fsm_output[1]);
      D_1_5_sva <= MUX_s_1_2_2((key_rsci_idat[51]), D_1_5_sva_mx1, fsm_output[1]);
      D_1_6_sva <= MUX_s_1_2_2((key_rsci_idat[43]), D_1_6_sva_mx1, fsm_output[1]);
      D_1_7_sva <= MUX_s_1_2_2((key_rsci_idat[35]), D_1_7_sva_mx1, fsm_output[1]);
      D_1_8_sva <= MUX_s_1_2_2((key_rsci_idat[27]), D_1_8_sva_mx1, fsm_output[1]);
      D_1_9_sva <= MUX_s_1_2_2((key_rsci_idat[19]), D_1_9_sva_mx1, fsm_output[1]);
      D_1_10_sva <= MUX_s_1_2_2((key_rsci_idat[11]), D_1_10_sva_mx1, fsm_output[1]);
      D_1_11_sva <= MUX_s_1_2_2((key_rsci_idat[3]), D_1_11_sva_mx1, fsm_output[1]);
      D_1_12_sva <= MUX_s_1_2_2((key_rsci_idat[58]), D_1_12_sva_mx1, fsm_output[1]);
      D_1_13_sva <= MUX_s_1_2_2((key_rsci_idat[50]), D_mux_31_nl, fsm_output[1]);
      D_1_14_sva <= MUX_s_1_2_2((key_rsci_idat[42]), D_1_14_sva_mx1, fsm_output[1]);
      D_1_15_sva <= MUX_s_1_2_2((key_rsci_idat[34]), D_1_15_sva_mx1, fsm_output[1]);
      D_1_16_sva <= MUX_s_1_2_2((key_rsci_idat[26]), D_1_16_sva_mx1, fsm_output[1]);
      D_1_17_sva <= MUX_s_1_2_2((key_rsci_idat[18]), D_1_17_sva_mx1, fsm_output[1]);
      D_1_18_sva <= MUX_s_1_2_2((key_rsci_idat[10]), D_mux_41_nl, fsm_output[1]);
      D_1_19_sva <= MUX_s_1_2_2((key_rsci_idat[2]), D_1_19_sva_mx1, fsm_output[1]);
      D_1_20_sva <= MUX_s_1_2_2((key_rsci_idat[57]), D_1_20_sva_mx1, fsm_output[1]);
      D_1_21_sva <= MUX_s_1_2_2((key_rsci_idat[49]), D_mux_47_nl, fsm_output[1]);
      D_1_22_sva <= MUX_s_1_2_2((key_rsci_idat[41]), D_1_22_sva_mx1, fsm_output[1]);
      D_1_23_sva <= MUX_s_1_2_2((key_rsci_idat[33]), D_1_23_sva_mx1, fsm_output[1]);
      D_1_24_sva <= MUX_s_1_2_2((key_rsci_idat[25]), D_1_24_sva_mx1, fsm_output[1]);
      D_1_25_sva <= MUX_s_1_2_2((key_rsci_idat[17]), D_1_25_sva_mx1, fsm_output[1]);
      C_1_26_sva <= MUX_s_1_2_2((key_rsci_idat[15]), C_1_26_sva_mx1, fsm_output[1]);
      C_1_27_sva <= MUX_s_1_2_2((key_rsci_idat[7]), C_1_27_sva_mx1, fsm_output[1]);
      C_1_0_sva <= MUX_s_1_2_2((key_rsci_idat[28]), C_1_0_sva_mx1, fsm_output[1]);
      C_1_1_sva <= MUX_s_1_2_2((key_rsci_idat[20]), C_1_1_sva_mx1, fsm_output[1]);
      C_1_2_sva <= MUX_s_1_2_2((key_rsci_idat[12]), C_1_2_sva_mx1, fsm_output[1]);
      C_1_3_sva <= MUX_s_1_2_2((key_rsci_idat[4]), C_mux_11_nl, fsm_output[1]);
      C_1_4_sva <= MUX_s_1_2_2((key_rsci_idat[61]), C_1_4_sva_mx1, fsm_output[1]);
      C_1_5_sva <= MUX_s_1_2_2((key_rsci_idat[53]), C_1_5_sva_mx1, fsm_output[1]);
      C_1_6_sva <= MUX_s_1_2_2((key_rsci_idat[45]), C_mux_17_nl, fsm_output[1]);
      C_1_7_sva <= MUX_s_1_2_2((key_rsci_idat[37]), C_1_7_sva_mx1, fsm_output[1]);
      C_1_8_sva <= MUX_s_1_2_2((key_rsci_idat[29]), C_1_8_sva_mx1, fsm_output[1]);
      C_1_9_sva <= MUX_s_1_2_2((key_rsci_idat[21]), C_1_9_sva_mx1, fsm_output[1]);
      C_1_10_sva <= MUX_s_1_2_2((key_rsci_idat[13]), C_mux_25_nl, fsm_output[1]);
      C_1_11_sva <= MUX_s_1_2_2((key_rsci_idat[5]), C_1_11_sva_mx1, fsm_output[1]);
      C_1_12_sva <= MUX_s_1_2_2((key_rsci_idat[62]), C_1_12_sva_mx1, fsm_output[1]);
      C_1_13_sva <= MUX_s_1_2_2((key_rsci_idat[54]), C_1_13_sva_mx1, fsm_output[1]);
      C_1_14_sva <= MUX_s_1_2_2((key_rsci_idat[46]), C_1_14_sva_mx1, fsm_output[1]);
      C_1_15_sva <= MUX_s_1_2_2((key_rsci_idat[38]), C_1_15_sva_mx1, fsm_output[1]);
      C_1_16_sva <= MUX_s_1_2_2((key_rsci_idat[30]), C_1_16_sva_mx1, fsm_output[1]);
      C_1_17_sva <= MUX_s_1_2_2((key_rsci_idat[22]), C_1_17_sva_mx1, fsm_output[1]);
      C_1_18_sva <= MUX_s_1_2_2((key_rsci_idat[14]), C_1_18_sva_mx1, fsm_output[1]);
      C_1_19_sva <= MUX_s_1_2_2((key_rsci_idat[6]), C_mux_43_nl, fsm_output[1]);
      C_1_20_sva <= MUX_s_1_2_2((key_rsci_idat[63]), C_1_20_sva_mx1, fsm_output[1]);
      C_1_21_sva <= MUX_s_1_2_2((key_rsci_idat[55]), C_1_21_sva_mx1, fsm_output[1]);
      C_1_22_sva <= MUX_s_1_2_2((key_rsci_idat[47]), C_1_22_sva_mx1, fsm_output[1]);
      C_1_23_sva <= MUX_s_1_2_2((key_rsci_idat[39]), C_1_23_sva_mx1, fsm_output[1]);
      C_1_24_sva <= MUX_s_1_2_2((key_rsci_idat[31]), C_1_24_sva_mx1, fsm_output[1]);
      C_1_25_sva <= MUX_s_1_2_2((key_rsci_idat[23]), C_1_25_sva_mx1, fsm_output[1]);
      reg_return_rsc_triosy_obj_ld_cse <= (i_3_4_0_sva_2[4]) & (fsm_output[1]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_0 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_0 <= R_7_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_1 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_1 <= R_7_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_2 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_2 <= R_15_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_3 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_3 <= R_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_4 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_4 <= R_23_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_5 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_5 <= R_23_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_6 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_6 <= R_31_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_7 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_7 <= R_31_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_8 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_8 <= R_6_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_9 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_9 <= R_6_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_10 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_10 <= R_14_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_11 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_11 <= R_14_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_12 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_12 <= R_22_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_13 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_13 <= R_22_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_14 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_14 <= R_30_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_15 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_15 <= R_30_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_16 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_16 <= R_5_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_17 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_17 <= R_5_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_18 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_18 <= R_13_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_19 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_19 <= R_13_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_20 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_20 <= R_21_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_21 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_21 <= R_21_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_22 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_22 <= R_29_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_23 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_23 <= R_29_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_24 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_24 <= R_4_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_25 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_25 <= R_4_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_26 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_26 <= R_12_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_27 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_27 <= R_12_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_28 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_28 <= R_20_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_29 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_29 <= R_20_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_30 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_30 <= R_28_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_31 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_31 <= R_28_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_32 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_32 <= R_3_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_33 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_33 <= R_3_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_34 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_34 <= R_11_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_35 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_35 <= R_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_36 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_36 <= R_19_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_37 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_37 <= R_19_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_38 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_38 <= R_27_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_39 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_39 <= R_27_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_40 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_40 <= R_2_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_41 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_41 <= R_2_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_42 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_42 <= R_10_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_43 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_43 <= R_10_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_44 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_44 <= R_18_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_45 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_45 <= R_18_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_46 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_46 <= R_26_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_47 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_47 <= R_26_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_48 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_48 <= R_1_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_49 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_49 <= R_1_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_50 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_50 <= R_9_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_51 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_51 <= R_9_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_52 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_52 <= R_17_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_53 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_53 <= R_17_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_54 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_54 <= R_25_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_55 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_55 <= R_25_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_56 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_56 <= R_0_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_57 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_57 <= R_0_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_58 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_58 <= R_8_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_59 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_59 <= R_8_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_60 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_60 <= R_16_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_61 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_61 <= R_16_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_62 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_62 <= R_24_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsci_idat_63 <= 1'b0;
    end
    else if ( ~ or_tmp_121 ) begin
      return_rsci_idat_63 <= R_24_sva;
    end
  end
  assign D_mux_9_nl = MUX_s_1_2_2(D_1_1_sva, D_1_0_sva, not_tmp_1);
  assign D_mux_31_nl = MUX_s_1_2_2(D_1_12_sva, D_1_11_sva, not_tmp_1);
  assign D_mux_41_nl = MUX_s_1_2_2(D_1_17_sva, D_1_16_sva, not_tmp_1);
  assign D_mux_47_nl = MUX_s_1_2_2(D_1_20_sva, D_1_19_sva, not_tmp_1);
  assign C_mux_11_nl = MUX_s_1_2_2(C_1_2_sva, C_1_1_sva, not_tmp_1);
  assign C_mux_17_nl = MUX_s_1_2_2(C_1_5_sva, C_1_4_sva, not_tmp_1);
  assign C_mux_25_nl = MUX_s_1_2_2(C_1_9_sva, C_1_8_sva, not_tmp_1);
  assign C_mux_43_nl = MUX_s_1_2_2(C_1_18_sva, C_1_17_sva, not_tmp_1);

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    des_check
// ------------------------------------------------------------------


module des_check (
  clk, rst, input_rsc_dat, input_rsc_triosy_lz, key_rsc_dat, key_rsc_triosy_lz, return_rsc_dat,
      return_rsc_triosy_lz
);
  input clk;
  input rst;
  input [63:0] input_rsc_dat;
  output input_rsc_triosy_lz;
  input [63:0] key_rsc_dat;
  output key_rsc_triosy_lz;
  output [63:0] return_rsc_dat;
  output return_rsc_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  des_check_core des_check_core_inst (
      .clk(clk),
      .rst(rst),
      .input_rsc_dat(input_rsc_dat),
      .input_rsc_triosy_lz(input_rsc_triosy_lz),
      .key_rsc_dat(key_rsc_dat),
      .key_rsc_triosy_lz(key_rsc_triosy_lz),
      .return_rsc_dat(return_rsc_dat),
      .return_rsc_triosy_lz(return_rsc_triosy_lz)
    );
endmodule



